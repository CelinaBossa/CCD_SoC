magic
tech sky130A
magscale 1 2
timestamp 1723064828
<< pwell >>
rect -9679 -358 9679 358
<< mvnmos >>
rect -9451 -100 -9351 100
rect -9293 -100 -9193 100
rect -9135 -100 -9035 100
rect -8977 -100 -8877 100
rect -8819 -100 -8719 100
rect -8661 -100 -8561 100
rect -8503 -100 -8403 100
rect -8345 -100 -8245 100
rect -8187 -100 -8087 100
rect -8029 -100 -7929 100
rect -7871 -100 -7771 100
rect -7713 -100 -7613 100
rect -7555 -100 -7455 100
rect -7397 -100 -7297 100
rect -7239 -100 -7139 100
rect -7081 -100 -6981 100
rect -6923 -100 -6823 100
rect -6765 -100 -6665 100
rect -6607 -100 -6507 100
rect -6449 -100 -6349 100
rect -6291 -100 -6191 100
rect -6133 -100 -6033 100
rect -5975 -100 -5875 100
rect -5817 -100 -5717 100
rect -5659 -100 -5559 100
rect -5501 -100 -5401 100
rect -5343 -100 -5243 100
rect -5185 -100 -5085 100
rect -5027 -100 -4927 100
rect -4869 -100 -4769 100
rect -4711 -100 -4611 100
rect -4553 -100 -4453 100
rect -4395 -100 -4295 100
rect -4237 -100 -4137 100
rect -4079 -100 -3979 100
rect -3921 -100 -3821 100
rect -3763 -100 -3663 100
rect -3605 -100 -3505 100
rect -3447 -100 -3347 100
rect -3289 -100 -3189 100
rect -3131 -100 -3031 100
rect -2973 -100 -2873 100
rect -2815 -100 -2715 100
rect -2657 -100 -2557 100
rect -2499 -100 -2399 100
rect -2341 -100 -2241 100
rect -2183 -100 -2083 100
rect -2025 -100 -1925 100
rect -1867 -100 -1767 100
rect -1709 -100 -1609 100
rect -1551 -100 -1451 100
rect -1393 -100 -1293 100
rect -1235 -100 -1135 100
rect -1077 -100 -977 100
rect -919 -100 -819 100
rect -761 -100 -661 100
rect -603 -100 -503 100
rect -445 -100 -345 100
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
rect 345 -100 445 100
rect 503 -100 603 100
rect 661 -100 761 100
rect 819 -100 919 100
rect 977 -100 1077 100
rect 1135 -100 1235 100
rect 1293 -100 1393 100
rect 1451 -100 1551 100
rect 1609 -100 1709 100
rect 1767 -100 1867 100
rect 1925 -100 2025 100
rect 2083 -100 2183 100
rect 2241 -100 2341 100
rect 2399 -100 2499 100
rect 2557 -100 2657 100
rect 2715 -100 2815 100
rect 2873 -100 2973 100
rect 3031 -100 3131 100
rect 3189 -100 3289 100
rect 3347 -100 3447 100
rect 3505 -100 3605 100
rect 3663 -100 3763 100
rect 3821 -100 3921 100
rect 3979 -100 4079 100
rect 4137 -100 4237 100
rect 4295 -100 4395 100
rect 4453 -100 4553 100
rect 4611 -100 4711 100
rect 4769 -100 4869 100
rect 4927 -100 5027 100
rect 5085 -100 5185 100
rect 5243 -100 5343 100
rect 5401 -100 5501 100
rect 5559 -100 5659 100
rect 5717 -100 5817 100
rect 5875 -100 5975 100
rect 6033 -100 6133 100
rect 6191 -100 6291 100
rect 6349 -100 6449 100
rect 6507 -100 6607 100
rect 6665 -100 6765 100
rect 6823 -100 6923 100
rect 6981 -100 7081 100
rect 7139 -100 7239 100
rect 7297 -100 7397 100
rect 7455 -100 7555 100
rect 7613 -100 7713 100
rect 7771 -100 7871 100
rect 7929 -100 8029 100
rect 8087 -100 8187 100
rect 8245 -100 8345 100
rect 8403 -100 8503 100
rect 8561 -100 8661 100
rect 8719 -100 8819 100
rect 8877 -100 8977 100
rect 9035 -100 9135 100
rect 9193 -100 9293 100
rect 9351 -100 9451 100
<< mvndiff >>
rect -9509 88 -9451 100
rect -9509 -88 -9497 88
rect -9463 -88 -9451 88
rect -9509 -100 -9451 -88
rect -9351 88 -9293 100
rect -9351 -88 -9339 88
rect -9305 -88 -9293 88
rect -9351 -100 -9293 -88
rect -9193 88 -9135 100
rect -9193 -88 -9181 88
rect -9147 -88 -9135 88
rect -9193 -100 -9135 -88
rect -9035 88 -8977 100
rect -9035 -88 -9023 88
rect -8989 -88 -8977 88
rect -9035 -100 -8977 -88
rect -8877 88 -8819 100
rect -8877 -88 -8865 88
rect -8831 -88 -8819 88
rect -8877 -100 -8819 -88
rect -8719 88 -8661 100
rect -8719 -88 -8707 88
rect -8673 -88 -8661 88
rect -8719 -100 -8661 -88
rect -8561 88 -8503 100
rect -8561 -88 -8549 88
rect -8515 -88 -8503 88
rect -8561 -100 -8503 -88
rect -8403 88 -8345 100
rect -8403 -88 -8391 88
rect -8357 -88 -8345 88
rect -8403 -100 -8345 -88
rect -8245 88 -8187 100
rect -8245 -88 -8233 88
rect -8199 -88 -8187 88
rect -8245 -100 -8187 -88
rect -8087 88 -8029 100
rect -8087 -88 -8075 88
rect -8041 -88 -8029 88
rect -8087 -100 -8029 -88
rect -7929 88 -7871 100
rect -7929 -88 -7917 88
rect -7883 -88 -7871 88
rect -7929 -100 -7871 -88
rect -7771 88 -7713 100
rect -7771 -88 -7759 88
rect -7725 -88 -7713 88
rect -7771 -100 -7713 -88
rect -7613 88 -7555 100
rect -7613 -88 -7601 88
rect -7567 -88 -7555 88
rect -7613 -100 -7555 -88
rect -7455 88 -7397 100
rect -7455 -88 -7443 88
rect -7409 -88 -7397 88
rect -7455 -100 -7397 -88
rect -7297 88 -7239 100
rect -7297 -88 -7285 88
rect -7251 -88 -7239 88
rect -7297 -100 -7239 -88
rect -7139 88 -7081 100
rect -7139 -88 -7127 88
rect -7093 -88 -7081 88
rect -7139 -100 -7081 -88
rect -6981 88 -6923 100
rect -6981 -88 -6969 88
rect -6935 -88 -6923 88
rect -6981 -100 -6923 -88
rect -6823 88 -6765 100
rect -6823 -88 -6811 88
rect -6777 -88 -6765 88
rect -6823 -100 -6765 -88
rect -6665 88 -6607 100
rect -6665 -88 -6653 88
rect -6619 -88 -6607 88
rect -6665 -100 -6607 -88
rect -6507 88 -6449 100
rect -6507 -88 -6495 88
rect -6461 -88 -6449 88
rect -6507 -100 -6449 -88
rect -6349 88 -6291 100
rect -6349 -88 -6337 88
rect -6303 -88 -6291 88
rect -6349 -100 -6291 -88
rect -6191 88 -6133 100
rect -6191 -88 -6179 88
rect -6145 -88 -6133 88
rect -6191 -100 -6133 -88
rect -6033 88 -5975 100
rect -6033 -88 -6021 88
rect -5987 -88 -5975 88
rect -6033 -100 -5975 -88
rect -5875 88 -5817 100
rect -5875 -88 -5863 88
rect -5829 -88 -5817 88
rect -5875 -100 -5817 -88
rect -5717 88 -5659 100
rect -5717 -88 -5705 88
rect -5671 -88 -5659 88
rect -5717 -100 -5659 -88
rect -5559 88 -5501 100
rect -5559 -88 -5547 88
rect -5513 -88 -5501 88
rect -5559 -100 -5501 -88
rect -5401 88 -5343 100
rect -5401 -88 -5389 88
rect -5355 -88 -5343 88
rect -5401 -100 -5343 -88
rect -5243 88 -5185 100
rect -5243 -88 -5231 88
rect -5197 -88 -5185 88
rect -5243 -100 -5185 -88
rect -5085 88 -5027 100
rect -5085 -88 -5073 88
rect -5039 -88 -5027 88
rect -5085 -100 -5027 -88
rect -4927 88 -4869 100
rect -4927 -88 -4915 88
rect -4881 -88 -4869 88
rect -4927 -100 -4869 -88
rect -4769 88 -4711 100
rect -4769 -88 -4757 88
rect -4723 -88 -4711 88
rect -4769 -100 -4711 -88
rect -4611 88 -4553 100
rect -4611 -88 -4599 88
rect -4565 -88 -4553 88
rect -4611 -100 -4553 -88
rect -4453 88 -4395 100
rect -4453 -88 -4441 88
rect -4407 -88 -4395 88
rect -4453 -100 -4395 -88
rect -4295 88 -4237 100
rect -4295 -88 -4283 88
rect -4249 -88 -4237 88
rect -4295 -100 -4237 -88
rect -4137 88 -4079 100
rect -4137 -88 -4125 88
rect -4091 -88 -4079 88
rect -4137 -100 -4079 -88
rect -3979 88 -3921 100
rect -3979 -88 -3967 88
rect -3933 -88 -3921 88
rect -3979 -100 -3921 -88
rect -3821 88 -3763 100
rect -3821 -88 -3809 88
rect -3775 -88 -3763 88
rect -3821 -100 -3763 -88
rect -3663 88 -3605 100
rect -3663 -88 -3651 88
rect -3617 -88 -3605 88
rect -3663 -100 -3605 -88
rect -3505 88 -3447 100
rect -3505 -88 -3493 88
rect -3459 -88 -3447 88
rect -3505 -100 -3447 -88
rect -3347 88 -3289 100
rect -3347 -88 -3335 88
rect -3301 -88 -3289 88
rect -3347 -100 -3289 -88
rect -3189 88 -3131 100
rect -3189 -88 -3177 88
rect -3143 -88 -3131 88
rect -3189 -100 -3131 -88
rect -3031 88 -2973 100
rect -3031 -88 -3019 88
rect -2985 -88 -2973 88
rect -3031 -100 -2973 -88
rect -2873 88 -2815 100
rect -2873 -88 -2861 88
rect -2827 -88 -2815 88
rect -2873 -100 -2815 -88
rect -2715 88 -2657 100
rect -2715 -88 -2703 88
rect -2669 -88 -2657 88
rect -2715 -100 -2657 -88
rect -2557 88 -2499 100
rect -2557 -88 -2545 88
rect -2511 -88 -2499 88
rect -2557 -100 -2499 -88
rect -2399 88 -2341 100
rect -2399 -88 -2387 88
rect -2353 -88 -2341 88
rect -2399 -100 -2341 -88
rect -2241 88 -2183 100
rect -2241 -88 -2229 88
rect -2195 -88 -2183 88
rect -2241 -100 -2183 -88
rect -2083 88 -2025 100
rect -2083 -88 -2071 88
rect -2037 -88 -2025 88
rect -2083 -100 -2025 -88
rect -1925 88 -1867 100
rect -1925 -88 -1913 88
rect -1879 -88 -1867 88
rect -1925 -100 -1867 -88
rect -1767 88 -1709 100
rect -1767 -88 -1755 88
rect -1721 -88 -1709 88
rect -1767 -100 -1709 -88
rect -1609 88 -1551 100
rect -1609 -88 -1597 88
rect -1563 -88 -1551 88
rect -1609 -100 -1551 -88
rect -1451 88 -1393 100
rect -1451 -88 -1439 88
rect -1405 -88 -1393 88
rect -1451 -100 -1393 -88
rect -1293 88 -1235 100
rect -1293 -88 -1281 88
rect -1247 -88 -1235 88
rect -1293 -100 -1235 -88
rect -1135 88 -1077 100
rect -1135 -88 -1123 88
rect -1089 -88 -1077 88
rect -1135 -100 -1077 -88
rect -977 88 -919 100
rect -977 -88 -965 88
rect -931 -88 -919 88
rect -977 -100 -919 -88
rect -819 88 -761 100
rect -819 -88 -807 88
rect -773 -88 -761 88
rect -819 -100 -761 -88
rect -661 88 -603 100
rect -661 -88 -649 88
rect -615 -88 -603 88
rect -661 -100 -603 -88
rect -503 88 -445 100
rect -503 -88 -491 88
rect -457 -88 -445 88
rect -503 -100 -445 -88
rect -345 88 -287 100
rect -345 -88 -333 88
rect -299 -88 -287 88
rect -345 -100 -287 -88
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
rect 287 88 345 100
rect 287 -88 299 88
rect 333 -88 345 88
rect 287 -100 345 -88
rect 445 88 503 100
rect 445 -88 457 88
rect 491 -88 503 88
rect 445 -100 503 -88
rect 603 88 661 100
rect 603 -88 615 88
rect 649 -88 661 88
rect 603 -100 661 -88
rect 761 88 819 100
rect 761 -88 773 88
rect 807 -88 819 88
rect 761 -100 819 -88
rect 919 88 977 100
rect 919 -88 931 88
rect 965 -88 977 88
rect 919 -100 977 -88
rect 1077 88 1135 100
rect 1077 -88 1089 88
rect 1123 -88 1135 88
rect 1077 -100 1135 -88
rect 1235 88 1293 100
rect 1235 -88 1247 88
rect 1281 -88 1293 88
rect 1235 -100 1293 -88
rect 1393 88 1451 100
rect 1393 -88 1405 88
rect 1439 -88 1451 88
rect 1393 -100 1451 -88
rect 1551 88 1609 100
rect 1551 -88 1563 88
rect 1597 -88 1609 88
rect 1551 -100 1609 -88
rect 1709 88 1767 100
rect 1709 -88 1721 88
rect 1755 -88 1767 88
rect 1709 -100 1767 -88
rect 1867 88 1925 100
rect 1867 -88 1879 88
rect 1913 -88 1925 88
rect 1867 -100 1925 -88
rect 2025 88 2083 100
rect 2025 -88 2037 88
rect 2071 -88 2083 88
rect 2025 -100 2083 -88
rect 2183 88 2241 100
rect 2183 -88 2195 88
rect 2229 -88 2241 88
rect 2183 -100 2241 -88
rect 2341 88 2399 100
rect 2341 -88 2353 88
rect 2387 -88 2399 88
rect 2341 -100 2399 -88
rect 2499 88 2557 100
rect 2499 -88 2511 88
rect 2545 -88 2557 88
rect 2499 -100 2557 -88
rect 2657 88 2715 100
rect 2657 -88 2669 88
rect 2703 -88 2715 88
rect 2657 -100 2715 -88
rect 2815 88 2873 100
rect 2815 -88 2827 88
rect 2861 -88 2873 88
rect 2815 -100 2873 -88
rect 2973 88 3031 100
rect 2973 -88 2985 88
rect 3019 -88 3031 88
rect 2973 -100 3031 -88
rect 3131 88 3189 100
rect 3131 -88 3143 88
rect 3177 -88 3189 88
rect 3131 -100 3189 -88
rect 3289 88 3347 100
rect 3289 -88 3301 88
rect 3335 -88 3347 88
rect 3289 -100 3347 -88
rect 3447 88 3505 100
rect 3447 -88 3459 88
rect 3493 -88 3505 88
rect 3447 -100 3505 -88
rect 3605 88 3663 100
rect 3605 -88 3617 88
rect 3651 -88 3663 88
rect 3605 -100 3663 -88
rect 3763 88 3821 100
rect 3763 -88 3775 88
rect 3809 -88 3821 88
rect 3763 -100 3821 -88
rect 3921 88 3979 100
rect 3921 -88 3933 88
rect 3967 -88 3979 88
rect 3921 -100 3979 -88
rect 4079 88 4137 100
rect 4079 -88 4091 88
rect 4125 -88 4137 88
rect 4079 -100 4137 -88
rect 4237 88 4295 100
rect 4237 -88 4249 88
rect 4283 -88 4295 88
rect 4237 -100 4295 -88
rect 4395 88 4453 100
rect 4395 -88 4407 88
rect 4441 -88 4453 88
rect 4395 -100 4453 -88
rect 4553 88 4611 100
rect 4553 -88 4565 88
rect 4599 -88 4611 88
rect 4553 -100 4611 -88
rect 4711 88 4769 100
rect 4711 -88 4723 88
rect 4757 -88 4769 88
rect 4711 -100 4769 -88
rect 4869 88 4927 100
rect 4869 -88 4881 88
rect 4915 -88 4927 88
rect 4869 -100 4927 -88
rect 5027 88 5085 100
rect 5027 -88 5039 88
rect 5073 -88 5085 88
rect 5027 -100 5085 -88
rect 5185 88 5243 100
rect 5185 -88 5197 88
rect 5231 -88 5243 88
rect 5185 -100 5243 -88
rect 5343 88 5401 100
rect 5343 -88 5355 88
rect 5389 -88 5401 88
rect 5343 -100 5401 -88
rect 5501 88 5559 100
rect 5501 -88 5513 88
rect 5547 -88 5559 88
rect 5501 -100 5559 -88
rect 5659 88 5717 100
rect 5659 -88 5671 88
rect 5705 -88 5717 88
rect 5659 -100 5717 -88
rect 5817 88 5875 100
rect 5817 -88 5829 88
rect 5863 -88 5875 88
rect 5817 -100 5875 -88
rect 5975 88 6033 100
rect 5975 -88 5987 88
rect 6021 -88 6033 88
rect 5975 -100 6033 -88
rect 6133 88 6191 100
rect 6133 -88 6145 88
rect 6179 -88 6191 88
rect 6133 -100 6191 -88
rect 6291 88 6349 100
rect 6291 -88 6303 88
rect 6337 -88 6349 88
rect 6291 -100 6349 -88
rect 6449 88 6507 100
rect 6449 -88 6461 88
rect 6495 -88 6507 88
rect 6449 -100 6507 -88
rect 6607 88 6665 100
rect 6607 -88 6619 88
rect 6653 -88 6665 88
rect 6607 -100 6665 -88
rect 6765 88 6823 100
rect 6765 -88 6777 88
rect 6811 -88 6823 88
rect 6765 -100 6823 -88
rect 6923 88 6981 100
rect 6923 -88 6935 88
rect 6969 -88 6981 88
rect 6923 -100 6981 -88
rect 7081 88 7139 100
rect 7081 -88 7093 88
rect 7127 -88 7139 88
rect 7081 -100 7139 -88
rect 7239 88 7297 100
rect 7239 -88 7251 88
rect 7285 -88 7297 88
rect 7239 -100 7297 -88
rect 7397 88 7455 100
rect 7397 -88 7409 88
rect 7443 -88 7455 88
rect 7397 -100 7455 -88
rect 7555 88 7613 100
rect 7555 -88 7567 88
rect 7601 -88 7613 88
rect 7555 -100 7613 -88
rect 7713 88 7771 100
rect 7713 -88 7725 88
rect 7759 -88 7771 88
rect 7713 -100 7771 -88
rect 7871 88 7929 100
rect 7871 -88 7883 88
rect 7917 -88 7929 88
rect 7871 -100 7929 -88
rect 8029 88 8087 100
rect 8029 -88 8041 88
rect 8075 -88 8087 88
rect 8029 -100 8087 -88
rect 8187 88 8245 100
rect 8187 -88 8199 88
rect 8233 -88 8245 88
rect 8187 -100 8245 -88
rect 8345 88 8403 100
rect 8345 -88 8357 88
rect 8391 -88 8403 88
rect 8345 -100 8403 -88
rect 8503 88 8561 100
rect 8503 -88 8515 88
rect 8549 -88 8561 88
rect 8503 -100 8561 -88
rect 8661 88 8719 100
rect 8661 -88 8673 88
rect 8707 -88 8719 88
rect 8661 -100 8719 -88
rect 8819 88 8877 100
rect 8819 -88 8831 88
rect 8865 -88 8877 88
rect 8819 -100 8877 -88
rect 8977 88 9035 100
rect 8977 -88 8989 88
rect 9023 -88 9035 88
rect 8977 -100 9035 -88
rect 9135 88 9193 100
rect 9135 -88 9147 88
rect 9181 -88 9193 88
rect 9135 -100 9193 -88
rect 9293 88 9351 100
rect 9293 -88 9305 88
rect 9339 -88 9351 88
rect 9293 -100 9351 -88
rect 9451 88 9509 100
rect 9451 -88 9463 88
rect 9497 -88 9509 88
rect 9451 -100 9509 -88
<< mvndiffc >>
rect -9497 -88 -9463 88
rect -9339 -88 -9305 88
rect -9181 -88 -9147 88
rect -9023 -88 -8989 88
rect -8865 -88 -8831 88
rect -8707 -88 -8673 88
rect -8549 -88 -8515 88
rect -8391 -88 -8357 88
rect -8233 -88 -8199 88
rect -8075 -88 -8041 88
rect -7917 -88 -7883 88
rect -7759 -88 -7725 88
rect -7601 -88 -7567 88
rect -7443 -88 -7409 88
rect -7285 -88 -7251 88
rect -7127 -88 -7093 88
rect -6969 -88 -6935 88
rect -6811 -88 -6777 88
rect -6653 -88 -6619 88
rect -6495 -88 -6461 88
rect -6337 -88 -6303 88
rect -6179 -88 -6145 88
rect -6021 -88 -5987 88
rect -5863 -88 -5829 88
rect -5705 -88 -5671 88
rect -5547 -88 -5513 88
rect -5389 -88 -5355 88
rect -5231 -88 -5197 88
rect -5073 -88 -5039 88
rect -4915 -88 -4881 88
rect -4757 -88 -4723 88
rect -4599 -88 -4565 88
rect -4441 -88 -4407 88
rect -4283 -88 -4249 88
rect -4125 -88 -4091 88
rect -3967 -88 -3933 88
rect -3809 -88 -3775 88
rect -3651 -88 -3617 88
rect -3493 -88 -3459 88
rect -3335 -88 -3301 88
rect -3177 -88 -3143 88
rect -3019 -88 -2985 88
rect -2861 -88 -2827 88
rect -2703 -88 -2669 88
rect -2545 -88 -2511 88
rect -2387 -88 -2353 88
rect -2229 -88 -2195 88
rect -2071 -88 -2037 88
rect -1913 -88 -1879 88
rect -1755 -88 -1721 88
rect -1597 -88 -1563 88
rect -1439 -88 -1405 88
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
rect 1405 -88 1439 88
rect 1563 -88 1597 88
rect 1721 -88 1755 88
rect 1879 -88 1913 88
rect 2037 -88 2071 88
rect 2195 -88 2229 88
rect 2353 -88 2387 88
rect 2511 -88 2545 88
rect 2669 -88 2703 88
rect 2827 -88 2861 88
rect 2985 -88 3019 88
rect 3143 -88 3177 88
rect 3301 -88 3335 88
rect 3459 -88 3493 88
rect 3617 -88 3651 88
rect 3775 -88 3809 88
rect 3933 -88 3967 88
rect 4091 -88 4125 88
rect 4249 -88 4283 88
rect 4407 -88 4441 88
rect 4565 -88 4599 88
rect 4723 -88 4757 88
rect 4881 -88 4915 88
rect 5039 -88 5073 88
rect 5197 -88 5231 88
rect 5355 -88 5389 88
rect 5513 -88 5547 88
rect 5671 -88 5705 88
rect 5829 -88 5863 88
rect 5987 -88 6021 88
rect 6145 -88 6179 88
rect 6303 -88 6337 88
rect 6461 -88 6495 88
rect 6619 -88 6653 88
rect 6777 -88 6811 88
rect 6935 -88 6969 88
rect 7093 -88 7127 88
rect 7251 -88 7285 88
rect 7409 -88 7443 88
rect 7567 -88 7601 88
rect 7725 -88 7759 88
rect 7883 -88 7917 88
rect 8041 -88 8075 88
rect 8199 -88 8233 88
rect 8357 -88 8391 88
rect 8515 -88 8549 88
rect 8673 -88 8707 88
rect 8831 -88 8865 88
rect 8989 -88 9023 88
rect 9147 -88 9181 88
rect 9305 -88 9339 88
rect 9463 -88 9497 88
<< mvpsubdiff >>
rect -9643 310 9643 322
rect -9643 276 -9535 310
rect 9535 276 9643 310
rect -9643 264 9643 276
rect -9643 214 -9585 264
rect -9643 -214 -9631 214
rect -9597 -214 -9585 214
rect 9585 214 9643 264
rect -9643 -264 -9585 -214
rect 9585 -214 9597 214
rect 9631 -214 9643 214
rect 9585 -264 9643 -214
rect -9643 -276 9643 -264
rect -9643 -310 -9535 -276
rect 9535 -310 9643 -276
rect -9643 -322 9643 -310
<< mvpsubdiffcont >>
rect -9535 276 9535 310
rect -9631 -214 -9597 214
rect 9597 -214 9631 214
rect -9535 -310 9535 -276
<< poly >>
rect -9451 172 -9351 188
rect -9451 138 -9435 172
rect -9367 138 -9351 172
rect -9451 100 -9351 138
rect -9293 172 -9193 188
rect -9293 138 -9277 172
rect -9209 138 -9193 172
rect -9293 100 -9193 138
rect -9135 172 -9035 188
rect -9135 138 -9119 172
rect -9051 138 -9035 172
rect -9135 100 -9035 138
rect -8977 172 -8877 188
rect -8977 138 -8961 172
rect -8893 138 -8877 172
rect -8977 100 -8877 138
rect -8819 172 -8719 188
rect -8819 138 -8803 172
rect -8735 138 -8719 172
rect -8819 100 -8719 138
rect -8661 172 -8561 188
rect -8661 138 -8645 172
rect -8577 138 -8561 172
rect -8661 100 -8561 138
rect -8503 172 -8403 188
rect -8503 138 -8487 172
rect -8419 138 -8403 172
rect -8503 100 -8403 138
rect -8345 172 -8245 188
rect -8345 138 -8329 172
rect -8261 138 -8245 172
rect -8345 100 -8245 138
rect -8187 172 -8087 188
rect -8187 138 -8171 172
rect -8103 138 -8087 172
rect -8187 100 -8087 138
rect -8029 172 -7929 188
rect -8029 138 -8013 172
rect -7945 138 -7929 172
rect -8029 100 -7929 138
rect -7871 172 -7771 188
rect -7871 138 -7855 172
rect -7787 138 -7771 172
rect -7871 100 -7771 138
rect -7713 172 -7613 188
rect -7713 138 -7697 172
rect -7629 138 -7613 172
rect -7713 100 -7613 138
rect -7555 172 -7455 188
rect -7555 138 -7539 172
rect -7471 138 -7455 172
rect -7555 100 -7455 138
rect -7397 172 -7297 188
rect -7397 138 -7381 172
rect -7313 138 -7297 172
rect -7397 100 -7297 138
rect -7239 172 -7139 188
rect -7239 138 -7223 172
rect -7155 138 -7139 172
rect -7239 100 -7139 138
rect -7081 172 -6981 188
rect -7081 138 -7065 172
rect -6997 138 -6981 172
rect -7081 100 -6981 138
rect -6923 172 -6823 188
rect -6923 138 -6907 172
rect -6839 138 -6823 172
rect -6923 100 -6823 138
rect -6765 172 -6665 188
rect -6765 138 -6749 172
rect -6681 138 -6665 172
rect -6765 100 -6665 138
rect -6607 172 -6507 188
rect -6607 138 -6591 172
rect -6523 138 -6507 172
rect -6607 100 -6507 138
rect -6449 172 -6349 188
rect -6449 138 -6433 172
rect -6365 138 -6349 172
rect -6449 100 -6349 138
rect -6291 172 -6191 188
rect -6291 138 -6275 172
rect -6207 138 -6191 172
rect -6291 100 -6191 138
rect -6133 172 -6033 188
rect -6133 138 -6117 172
rect -6049 138 -6033 172
rect -6133 100 -6033 138
rect -5975 172 -5875 188
rect -5975 138 -5959 172
rect -5891 138 -5875 172
rect -5975 100 -5875 138
rect -5817 172 -5717 188
rect -5817 138 -5801 172
rect -5733 138 -5717 172
rect -5817 100 -5717 138
rect -5659 172 -5559 188
rect -5659 138 -5643 172
rect -5575 138 -5559 172
rect -5659 100 -5559 138
rect -5501 172 -5401 188
rect -5501 138 -5485 172
rect -5417 138 -5401 172
rect -5501 100 -5401 138
rect -5343 172 -5243 188
rect -5343 138 -5327 172
rect -5259 138 -5243 172
rect -5343 100 -5243 138
rect -5185 172 -5085 188
rect -5185 138 -5169 172
rect -5101 138 -5085 172
rect -5185 100 -5085 138
rect -5027 172 -4927 188
rect -5027 138 -5011 172
rect -4943 138 -4927 172
rect -5027 100 -4927 138
rect -4869 172 -4769 188
rect -4869 138 -4853 172
rect -4785 138 -4769 172
rect -4869 100 -4769 138
rect -4711 172 -4611 188
rect -4711 138 -4695 172
rect -4627 138 -4611 172
rect -4711 100 -4611 138
rect -4553 172 -4453 188
rect -4553 138 -4537 172
rect -4469 138 -4453 172
rect -4553 100 -4453 138
rect -4395 172 -4295 188
rect -4395 138 -4379 172
rect -4311 138 -4295 172
rect -4395 100 -4295 138
rect -4237 172 -4137 188
rect -4237 138 -4221 172
rect -4153 138 -4137 172
rect -4237 100 -4137 138
rect -4079 172 -3979 188
rect -4079 138 -4063 172
rect -3995 138 -3979 172
rect -4079 100 -3979 138
rect -3921 172 -3821 188
rect -3921 138 -3905 172
rect -3837 138 -3821 172
rect -3921 100 -3821 138
rect -3763 172 -3663 188
rect -3763 138 -3747 172
rect -3679 138 -3663 172
rect -3763 100 -3663 138
rect -3605 172 -3505 188
rect -3605 138 -3589 172
rect -3521 138 -3505 172
rect -3605 100 -3505 138
rect -3447 172 -3347 188
rect -3447 138 -3431 172
rect -3363 138 -3347 172
rect -3447 100 -3347 138
rect -3289 172 -3189 188
rect -3289 138 -3273 172
rect -3205 138 -3189 172
rect -3289 100 -3189 138
rect -3131 172 -3031 188
rect -3131 138 -3115 172
rect -3047 138 -3031 172
rect -3131 100 -3031 138
rect -2973 172 -2873 188
rect -2973 138 -2957 172
rect -2889 138 -2873 172
rect -2973 100 -2873 138
rect -2815 172 -2715 188
rect -2815 138 -2799 172
rect -2731 138 -2715 172
rect -2815 100 -2715 138
rect -2657 172 -2557 188
rect -2657 138 -2641 172
rect -2573 138 -2557 172
rect -2657 100 -2557 138
rect -2499 172 -2399 188
rect -2499 138 -2483 172
rect -2415 138 -2399 172
rect -2499 100 -2399 138
rect -2341 172 -2241 188
rect -2341 138 -2325 172
rect -2257 138 -2241 172
rect -2341 100 -2241 138
rect -2183 172 -2083 188
rect -2183 138 -2167 172
rect -2099 138 -2083 172
rect -2183 100 -2083 138
rect -2025 172 -1925 188
rect -2025 138 -2009 172
rect -1941 138 -1925 172
rect -2025 100 -1925 138
rect -1867 172 -1767 188
rect -1867 138 -1851 172
rect -1783 138 -1767 172
rect -1867 100 -1767 138
rect -1709 172 -1609 188
rect -1709 138 -1693 172
rect -1625 138 -1609 172
rect -1709 100 -1609 138
rect -1551 172 -1451 188
rect -1551 138 -1535 172
rect -1467 138 -1451 172
rect -1551 100 -1451 138
rect -1393 172 -1293 188
rect -1393 138 -1377 172
rect -1309 138 -1293 172
rect -1393 100 -1293 138
rect -1235 172 -1135 188
rect -1235 138 -1219 172
rect -1151 138 -1135 172
rect -1235 100 -1135 138
rect -1077 172 -977 188
rect -1077 138 -1061 172
rect -993 138 -977 172
rect -1077 100 -977 138
rect -919 172 -819 188
rect -919 138 -903 172
rect -835 138 -819 172
rect -919 100 -819 138
rect -761 172 -661 188
rect -761 138 -745 172
rect -677 138 -661 172
rect -761 100 -661 138
rect -603 172 -503 188
rect -603 138 -587 172
rect -519 138 -503 172
rect -603 100 -503 138
rect -445 172 -345 188
rect -445 138 -429 172
rect -361 138 -345 172
rect -445 100 -345 138
rect -287 172 -187 188
rect -287 138 -271 172
rect -203 138 -187 172
rect -287 100 -187 138
rect -129 172 -29 188
rect -129 138 -113 172
rect -45 138 -29 172
rect -129 100 -29 138
rect 29 172 129 188
rect 29 138 45 172
rect 113 138 129 172
rect 29 100 129 138
rect 187 172 287 188
rect 187 138 203 172
rect 271 138 287 172
rect 187 100 287 138
rect 345 172 445 188
rect 345 138 361 172
rect 429 138 445 172
rect 345 100 445 138
rect 503 172 603 188
rect 503 138 519 172
rect 587 138 603 172
rect 503 100 603 138
rect 661 172 761 188
rect 661 138 677 172
rect 745 138 761 172
rect 661 100 761 138
rect 819 172 919 188
rect 819 138 835 172
rect 903 138 919 172
rect 819 100 919 138
rect 977 172 1077 188
rect 977 138 993 172
rect 1061 138 1077 172
rect 977 100 1077 138
rect 1135 172 1235 188
rect 1135 138 1151 172
rect 1219 138 1235 172
rect 1135 100 1235 138
rect 1293 172 1393 188
rect 1293 138 1309 172
rect 1377 138 1393 172
rect 1293 100 1393 138
rect 1451 172 1551 188
rect 1451 138 1467 172
rect 1535 138 1551 172
rect 1451 100 1551 138
rect 1609 172 1709 188
rect 1609 138 1625 172
rect 1693 138 1709 172
rect 1609 100 1709 138
rect 1767 172 1867 188
rect 1767 138 1783 172
rect 1851 138 1867 172
rect 1767 100 1867 138
rect 1925 172 2025 188
rect 1925 138 1941 172
rect 2009 138 2025 172
rect 1925 100 2025 138
rect 2083 172 2183 188
rect 2083 138 2099 172
rect 2167 138 2183 172
rect 2083 100 2183 138
rect 2241 172 2341 188
rect 2241 138 2257 172
rect 2325 138 2341 172
rect 2241 100 2341 138
rect 2399 172 2499 188
rect 2399 138 2415 172
rect 2483 138 2499 172
rect 2399 100 2499 138
rect 2557 172 2657 188
rect 2557 138 2573 172
rect 2641 138 2657 172
rect 2557 100 2657 138
rect 2715 172 2815 188
rect 2715 138 2731 172
rect 2799 138 2815 172
rect 2715 100 2815 138
rect 2873 172 2973 188
rect 2873 138 2889 172
rect 2957 138 2973 172
rect 2873 100 2973 138
rect 3031 172 3131 188
rect 3031 138 3047 172
rect 3115 138 3131 172
rect 3031 100 3131 138
rect 3189 172 3289 188
rect 3189 138 3205 172
rect 3273 138 3289 172
rect 3189 100 3289 138
rect 3347 172 3447 188
rect 3347 138 3363 172
rect 3431 138 3447 172
rect 3347 100 3447 138
rect 3505 172 3605 188
rect 3505 138 3521 172
rect 3589 138 3605 172
rect 3505 100 3605 138
rect 3663 172 3763 188
rect 3663 138 3679 172
rect 3747 138 3763 172
rect 3663 100 3763 138
rect 3821 172 3921 188
rect 3821 138 3837 172
rect 3905 138 3921 172
rect 3821 100 3921 138
rect 3979 172 4079 188
rect 3979 138 3995 172
rect 4063 138 4079 172
rect 3979 100 4079 138
rect 4137 172 4237 188
rect 4137 138 4153 172
rect 4221 138 4237 172
rect 4137 100 4237 138
rect 4295 172 4395 188
rect 4295 138 4311 172
rect 4379 138 4395 172
rect 4295 100 4395 138
rect 4453 172 4553 188
rect 4453 138 4469 172
rect 4537 138 4553 172
rect 4453 100 4553 138
rect 4611 172 4711 188
rect 4611 138 4627 172
rect 4695 138 4711 172
rect 4611 100 4711 138
rect 4769 172 4869 188
rect 4769 138 4785 172
rect 4853 138 4869 172
rect 4769 100 4869 138
rect 4927 172 5027 188
rect 4927 138 4943 172
rect 5011 138 5027 172
rect 4927 100 5027 138
rect 5085 172 5185 188
rect 5085 138 5101 172
rect 5169 138 5185 172
rect 5085 100 5185 138
rect 5243 172 5343 188
rect 5243 138 5259 172
rect 5327 138 5343 172
rect 5243 100 5343 138
rect 5401 172 5501 188
rect 5401 138 5417 172
rect 5485 138 5501 172
rect 5401 100 5501 138
rect 5559 172 5659 188
rect 5559 138 5575 172
rect 5643 138 5659 172
rect 5559 100 5659 138
rect 5717 172 5817 188
rect 5717 138 5733 172
rect 5801 138 5817 172
rect 5717 100 5817 138
rect 5875 172 5975 188
rect 5875 138 5891 172
rect 5959 138 5975 172
rect 5875 100 5975 138
rect 6033 172 6133 188
rect 6033 138 6049 172
rect 6117 138 6133 172
rect 6033 100 6133 138
rect 6191 172 6291 188
rect 6191 138 6207 172
rect 6275 138 6291 172
rect 6191 100 6291 138
rect 6349 172 6449 188
rect 6349 138 6365 172
rect 6433 138 6449 172
rect 6349 100 6449 138
rect 6507 172 6607 188
rect 6507 138 6523 172
rect 6591 138 6607 172
rect 6507 100 6607 138
rect 6665 172 6765 188
rect 6665 138 6681 172
rect 6749 138 6765 172
rect 6665 100 6765 138
rect 6823 172 6923 188
rect 6823 138 6839 172
rect 6907 138 6923 172
rect 6823 100 6923 138
rect 6981 172 7081 188
rect 6981 138 6997 172
rect 7065 138 7081 172
rect 6981 100 7081 138
rect 7139 172 7239 188
rect 7139 138 7155 172
rect 7223 138 7239 172
rect 7139 100 7239 138
rect 7297 172 7397 188
rect 7297 138 7313 172
rect 7381 138 7397 172
rect 7297 100 7397 138
rect 7455 172 7555 188
rect 7455 138 7471 172
rect 7539 138 7555 172
rect 7455 100 7555 138
rect 7613 172 7713 188
rect 7613 138 7629 172
rect 7697 138 7713 172
rect 7613 100 7713 138
rect 7771 172 7871 188
rect 7771 138 7787 172
rect 7855 138 7871 172
rect 7771 100 7871 138
rect 7929 172 8029 188
rect 7929 138 7945 172
rect 8013 138 8029 172
rect 7929 100 8029 138
rect 8087 172 8187 188
rect 8087 138 8103 172
rect 8171 138 8187 172
rect 8087 100 8187 138
rect 8245 172 8345 188
rect 8245 138 8261 172
rect 8329 138 8345 172
rect 8245 100 8345 138
rect 8403 172 8503 188
rect 8403 138 8419 172
rect 8487 138 8503 172
rect 8403 100 8503 138
rect 8561 172 8661 188
rect 8561 138 8577 172
rect 8645 138 8661 172
rect 8561 100 8661 138
rect 8719 172 8819 188
rect 8719 138 8735 172
rect 8803 138 8819 172
rect 8719 100 8819 138
rect 8877 172 8977 188
rect 8877 138 8893 172
rect 8961 138 8977 172
rect 8877 100 8977 138
rect 9035 172 9135 188
rect 9035 138 9051 172
rect 9119 138 9135 172
rect 9035 100 9135 138
rect 9193 172 9293 188
rect 9193 138 9209 172
rect 9277 138 9293 172
rect 9193 100 9293 138
rect 9351 172 9451 188
rect 9351 138 9367 172
rect 9435 138 9451 172
rect 9351 100 9451 138
rect -9451 -138 -9351 -100
rect -9451 -172 -9435 -138
rect -9367 -172 -9351 -138
rect -9451 -188 -9351 -172
rect -9293 -138 -9193 -100
rect -9293 -172 -9277 -138
rect -9209 -172 -9193 -138
rect -9293 -188 -9193 -172
rect -9135 -138 -9035 -100
rect -9135 -172 -9119 -138
rect -9051 -172 -9035 -138
rect -9135 -188 -9035 -172
rect -8977 -138 -8877 -100
rect -8977 -172 -8961 -138
rect -8893 -172 -8877 -138
rect -8977 -188 -8877 -172
rect -8819 -138 -8719 -100
rect -8819 -172 -8803 -138
rect -8735 -172 -8719 -138
rect -8819 -188 -8719 -172
rect -8661 -138 -8561 -100
rect -8661 -172 -8645 -138
rect -8577 -172 -8561 -138
rect -8661 -188 -8561 -172
rect -8503 -138 -8403 -100
rect -8503 -172 -8487 -138
rect -8419 -172 -8403 -138
rect -8503 -188 -8403 -172
rect -8345 -138 -8245 -100
rect -8345 -172 -8329 -138
rect -8261 -172 -8245 -138
rect -8345 -188 -8245 -172
rect -8187 -138 -8087 -100
rect -8187 -172 -8171 -138
rect -8103 -172 -8087 -138
rect -8187 -188 -8087 -172
rect -8029 -138 -7929 -100
rect -8029 -172 -8013 -138
rect -7945 -172 -7929 -138
rect -8029 -188 -7929 -172
rect -7871 -138 -7771 -100
rect -7871 -172 -7855 -138
rect -7787 -172 -7771 -138
rect -7871 -188 -7771 -172
rect -7713 -138 -7613 -100
rect -7713 -172 -7697 -138
rect -7629 -172 -7613 -138
rect -7713 -188 -7613 -172
rect -7555 -138 -7455 -100
rect -7555 -172 -7539 -138
rect -7471 -172 -7455 -138
rect -7555 -188 -7455 -172
rect -7397 -138 -7297 -100
rect -7397 -172 -7381 -138
rect -7313 -172 -7297 -138
rect -7397 -188 -7297 -172
rect -7239 -138 -7139 -100
rect -7239 -172 -7223 -138
rect -7155 -172 -7139 -138
rect -7239 -188 -7139 -172
rect -7081 -138 -6981 -100
rect -7081 -172 -7065 -138
rect -6997 -172 -6981 -138
rect -7081 -188 -6981 -172
rect -6923 -138 -6823 -100
rect -6923 -172 -6907 -138
rect -6839 -172 -6823 -138
rect -6923 -188 -6823 -172
rect -6765 -138 -6665 -100
rect -6765 -172 -6749 -138
rect -6681 -172 -6665 -138
rect -6765 -188 -6665 -172
rect -6607 -138 -6507 -100
rect -6607 -172 -6591 -138
rect -6523 -172 -6507 -138
rect -6607 -188 -6507 -172
rect -6449 -138 -6349 -100
rect -6449 -172 -6433 -138
rect -6365 -172 -6349 -138
rect -6449 -188 -6349 -172
rect -6291 -138 -6191 -100
rect -6291 -172 -6275 -138
rect -6207 -172 -6191 -138
rect -6291 -188 -6191 -172
rect -6133 -138 -6033 -100
rect -6133 -172 -6117 -138
rect -6049 -172 -6033 -138
rect -6133 -188 -6033 -172
rect -5975 -138 -5875 -100
rect -5975 -172 -5959 -138
rect -5891 -172 -5875 -138
rect -5975 -188 -5875 -172
rect -5817 -138 -5717 -100
rect -5817 -172 -5801 -138
rect -5733 -172 -5717 -138
rect -5817 -188 -5717 -172
rect -5659 -138 -5559 -100
rect -5659 -172 -5643 -138
rect -5575 -172 -5559 -138
rect -5659 -188 -5559 -172
rect -5501 -138 -5401 -100
rect -5501 -172 -5485 -138
rect -5417 -172 -5401 -138
rect -5501 -188 -5401 -172
rect -5343 -138 -5243 -100
rect -5343 -172 -5327 -138
rect -5259 -172 -5243 -138
rect -5343 -188 -5243 -172
rect -5185 -138 -5085 -100
rect -5185 -172 -5169 -138
rect -5101 -172 -5085 -138
rect -5185 -188 -5085 -172
rect -5027 -138 -4927 -100
rect -5027 -172 -5011 -138
rect -4943 -172 -4927 -138
rect -5027 -188 -4927 -172
rect -4869 -138 -4769 -100
rect -4869 -172 -4853 -138
rect -4785 -172 -4769 -138
rect -4869 -188 -4769 -172
rect -4711 -138 -4611 -100
rect -4711 -172 -4695 -138
rect -4627 -172 -4611 -138
rect -4711 -188 -4611 -172
rect -4553 -138 -4453 -100
rect -4553 -172 -4537 -138
rect -4469 -172 -4453 -138
rect -4553 -188 -4453 -172
rect -4395 -138 -4295 -100
rect -4395 -172 -4379 -138
rect -4311 -172 -4295 -138
rect -4395 -188 -4295 -172
rect -4237 -138 -4137 -100
rect -4237 -172 -4221 -138
rect -4153 -172 -4137 -138
rect -4237 -188 -4137 -172
rect -4079 -138 -3979 -100
rect -4079 -172 -4063 -138
rect -3995 -172 -3979 -138
rect -4079 -188 -3979 -172
rect -3921 -138 -3821 -100
rect -3921 -172 -3905 -138
rect -3837 -172 -3821 -138
rect -3921 -188 -3821 -172
rect -3763 -138 -3663 -100
rect -3763 -172 -3747 -138
rect -3679 -172 -3663 -138
rect -3763 -188 -3663 -172
rect -3605 -138 -3505 -100
rect -3605 -172 -3589 -138
rect -3521 -172 -3505 -138
rect -3605 -188 -3505 -172
rect -3447 -138 -3347 -100
rect -3447 -172 -3431 -138
rect -3363 -172 -3347 -138
rect -3447 -188 -3347 -172
rect -3289 -138 -3189 -100
rect -3289 -172 -3273 -138
rect -3205 -172 -3189 -138
rect -3289 -188 -3189 -172
rect -3131 -138 -3031 -100
rect -3131 -172 -3115 -138
rect -3047 -172 -3031 -138
rect -3131 -188 -3031 -172
rect -2973 -138 -2873 -100
rect -2973 -172 -2957 -138
rect -2889 -172 -2873 -138
rect -2973 -188 -2873 -172
rect -2815 -138 -2715 -100
rect -2815 -172 -2799 -138
rect -2731 -172 -2715 -138
rect -2815 -188 -2715 -172
rect -2657 -138 -2557 -100
rect -2657 -172 -2641 -138
rect -2573 -172 -2557 -138
rect -2657 -188 -2557 -172
rect -2499 -138 -2399 -100
rect -2499 -172 -2483 -138
rect -2415 -172 -2399 -138
rect -2499 -188 -2399 -172
rect -2341 -138 -2241 -100
rect -2341 -172 -2325 -138
rect -2257 -172 -2241 -138
rect -2341 -188 -2241 -172
rect -2183 -138 -2083 -100
rect -2183 -172 -2167 -138
rect -2099 -172 -2083 -138
rect -2183 -188 -2083 -172
rect -2025 -138 -1925 -100
rect -2025 -172 -2009 -138
rect -1941 -172 -1925 -138
rect -2025 -188 -1925 -172
rect -1867 -138 -1767 -100
rect -1867 -172 -1851 -138
rect -1783 -172 -1767 -138
rect -1867 -188 -1767 -172
rect -1709 -138 -1609 -100
rect -1709 -172 -1693 -138
rect -1625 -172 -1609 -138
rect -1709 -188 -1609 -172
rect -1551 -138 -1451 -100
rect -1551 -172 -1535 -138
rect -1467 -172 -1451 -138
rect -1551 -188 -1451 -172
rect -1393 -138 -1293 -100
rect -1393 -172 -1377 -138
rect -1309 -172 -1293 -138
rect -1393 -188 -1293 -172
rect -1235 -138 -1135 -100
rect -1235 -172 -1219 -138
rect -1151 -172 -1135 -138
rect -1235 -188 -1135 -172
rect -1077 -138 -977 -100
rect -1077 -172 -1061 -138
rect -993 -172 -977 -138
rect -1077 -188 -977 -172
rect -919 -138 -819 -100
rect -919 -172 -903 -138
rect -835 -172 -819 -138
rect -919 -188 -819 -172
rect -761 -138 -661 -100
rect -761 -172 -745 -138
rect -677 -172 -661 -138
rect -761 -188 -661 -172
rect -603 -138 -503 -100
rect -603 -172 -587 -138
rect -519 -172 -503 -138
rect -603 -188 -503 -172
rect -445 -138 -345 -100
rect -445 -172 -429 -138
rect -361 -172 -345 -138
rect -445 -188 -345 -172
rect -287 -138 -187 -100
rect -287 -172 -271 -138
rect -203 -172 -187 -138
rect -287 -188 -187 -172
rect -129 -138 -29 -100
rect -129 -172 -113 -138
rect -45 -172 -29 -138
rect -129 -188 -29 -172
rect 29 -138 129 -100
rect 29 -172 45 -138
rect 113 -172 129 -138
rect 29 -188 129 -172
rect 187 -138 287 -100
rect 187 -172 203 -138
rect 271 -172 287 -138
rect 187 -188 287 -172
rect 345 -138 445 -100
rect 345 -172 361 -138
rect 429 -172 445 -138
rect 345 -188 445 -172
rect 503 -138 603 -100
rect 503 -172 519 -138
rect 587 -172 603 -138
rect 503 -188 603 -172
rect 661 -138 761 -100
rect 661 -172 677 -138
rect 745 -172 761 -138
rect 661 -188 761 -172
rect 819 -138 919 -100
rect 819 -172 835 -138
rect 903 -172 919 -138
rect 819 -188 919 -172
rect 977 -138 1077 -100
rect 977 -172 993 -138
rect 1061 -172 1077 -138
rect 977 -188 1077 -172
rect 1135 -138 1235 -100
rect 1135 -172 1151 -138
rect 1219 -172 1235 -138
rect 1135 -188 1235 -172
rect 1293 -138 1393 -100
rect 1293 -172 1309 -138
rect 1377 -172 1393 -138
rect 1293 -188 1393 -172
rect 1451 -138 1551 -100
rect 1451 -172 1467 -138
rect 1535 -172 1551 -138
rect 1451 -188 1551 -172
rect 1609 -138 1709 -100
rect 1609 -172 1625 -138
rect 1693 -172 1709 -138
rect 1609 -188 1709 -172
rect 1767 -138 1867 -100
rect 1767 -172 1783 -138
rect 1851 -172 1867 -138
rect 1767 -188 1867 -172
rect 1925 -138 2025 -100
rect 1925 -172 1941 -138
rect 2009 -172 2025 -138
rect 1925 -188 2025 -172
rect 2083 -138 2183 -100
rect 2083 -172 2099 -138
rect 2167 -172 2183 -138
rect 2083 -188 2183 -172
rect 2241 -138 2341 -100
rect 2241 -172 2257 -138
rect 2325 -172 2341 -138
rect 2241 -188 2341 -172
rect 2399 -138 2499 -100
rect 2399 -172 2415 -138
rect 2483 -172 2499 -138
rect 2399 -188 2499 -172
rect 2557 -138 2657 -100
rect 2557 -172 2573 -138
rect 2641 -172 2657 -138
rect 2557 -188 2657 -172
rect 2715 -138 2815 -100
rect 2715 -172 2731 -138
rect 2799 -172 2815 -138
rect 2715 -188 2815 -172
rect 2873 -138 2973 -100
rect 2873 -172 2889 -138
rect 2957 -172 2973 -138
rect 2873 -188 2973 -172
rect 3031 -138 3131 -100
rect 3031 -172 3047 -138
rect 3115 -172 3131 -138
rect 3031 -188 3131 -172
rect 3189 -138 3289 -100
rect 3189 -172 3205 -138
rect 3273 -172 3289 -138
rect 3189 -188 3289 -172
rect 3347 -138 3447 -100
rect 3347 -172 3363 -138
rect 3431 -172 3447 -138
rect 3347 -188 3447 -172
rect 3505 -138 3605 -100
rect 3505 -172 3521 -138
rect 3589 -172 3605 -138
rect 3505 -188 3605 -172
rect 3663 -138 3763 -100
rect 3663 -172 3679 -138
rect 3747 -172 3763 -138
rect 3663 -188 3763 -172
rect 3821 -138 3921 -100
rect 3821 -172 3837 -138
rect 3905 -172 3921 -138
rect 3821 -188 3921 -172
rect 3979 -138 4079 -100
rect 3979 -172 3995 -138
rect 4063 -172 4079 -138
rect 3979 -188 4079 -172
rect 4137 -138 4237 -100
rect 4137 -172 4153 -138
rect 4221 -172 4237 -138
rect 4137 -188 4237 -172
rect 4295 -138 4395 -100
rect 4295 -172 4311 -138
rect 4379 -172 4395 -138
rect 4295 -188 4395 -172
rect 4453 -138 4553 -100
rect 4453 -172 4469 -138
rect 4537 -172 4553 -138
rect 4453 -188 4553 -172
rect 4611 -138 4711 -100
rect 4611 -172 4627 -138
rect 4695 -172 4711 -138
rect 4611 -188 4711 -172
rect 4769 -138 4869 -100
rect 4769 -172 4785 -138
rect 4853 -172 4869 -138
rect 4769 -188 4869 -172
rect 4927 -138 5027 -100
rect 4927 -172 4943 -138
rect 5011 -172 5027 -138
rect 4927 -188 5027 -172
rect 5085 -138 5185 -100
rect 5085 -172 5101 -138
rect 5169 -172 5185 -138
rect 5085 -188 5185 -172
rect 5243 -138 5343 -100
rect 5243 -172 5259 -138
rect 5327 -172 5343 -138
rect 5243 -188 5343 -172
rect 5401 -138 5501 -100
rect 5401 -172 5417 -138
rect 5485 -172 5501 -138
rect 5401 -188 5501 -172
rect 5559 -138 5659 -100
rect 5559 -172 5575 -138
rect 5643 -172 5659 -138
rect 5559 -188 5659 -172
rect 5717 -138 5817 -100
rect 5717 -172 5733 -138
rect 5801 -172 5817 -138
rect 5717 -188 5817 -172
rect 5875 -138 5975 -100
rect 5875 -172 5891 -138
rect 5959 -172 5975 -138
rect 5875 -188 5975 -172
rect 6033 -138 6133 -100
rect 6033 -172 6049 -138
rect 6117 -172 6133 -138
rect 6033 -188 6133 -172
rect 6191 -138 6291 -100
rect 6191 -172 6207 -138
rect 6275 -172 6291 -138
rect 6191 -188 6291 -172
rect 6349 -138 6449 -100
rect 6349 -172 6365 -138
rect 6433 -172 6449 -138
rect 6349 -188 6449 -172
rect 6507 -138 6607 -100
rect 6507 -172 6523 -138
rect 6591 -172 6607 -138
rect 6507 -188 6607 -172
rect 6665 -138 6765 -100
rect 6665 -172 6681 -138
rect 6749 -172 6765 -138
rect 6665 -188 6765 -172
rect 6823 -138 6923 -100
rect 6823 -172 6839 -138
rect 6907 -172 6923 -138
rect 6823 -188 6923 -172
rect 6981 -138 7081 -100
rect 6981 -172 6997 -138
rect 7065 -172 7081 -138
rect 6981 -188 7081 -172
rect 7139 -138 7239 -100
rect 7139 -172 7155 -138
rect 7223 -172 7239 -138
rect 7139 -188 7239 -172
rect 7297 -138 7397 -100
rect 7297 -172 7313 -138
rect 7381 -172 7397 -138
rect 7297 -188 7397 -172
rect 7455 -138 7555 -100
rect 7455 -172 7471 -138
rect 7539 -172 7555 -138
rect 7455 -188 7555 -172
rect 7613 -138 7713 -100
rect 7613 -172 7629 -138
rect 7697 -172 7713 -138
rect 7613 -188 7713 -172
rect 7771 -138 7871 -100
rect 7771 -172 7787 -138
rect 7855 -172 7871 -138
rect 7771 -188 7871 -172
rect 7929 -138 8029 -100
rect 7929 -172 7945 -138
rect 8013 -172 8029 -138
rect 7929 -188 8029 -172
rect 8087 -138 8187 -100
rect 8087 -172 8103 -138
rect 8171 -172 8187 -138
rect 8087 -188 8187 -172
rect 8245 -138 8345 -100
rect 8245 -172 8261 -138
rect 8329 -172 8345 -138
rect 8245 -188 8345 -172
rect 8403 -138 8503 -100
rect 8403 -172 8419 -138
rect 8487 -172 8503 -138
rect 8403 -188 8503 -172
rect 8561 -138 8661 -100
rect 8561 -172 8577 -138
rect 8645 -172 8661 -138
rect 8561 -188 8661 -172
rect 8719 -138 8819 -100
rect 8719 -172 8735 -138
rect 8803 -172 8819 -138
rect 8719 -188 8819 -172
rect 8877 -138 8977 -100
rect 8877 -172 8893 -138
rect 8961 -172 8977 -138
rect 8877 -188 8977 -172
rect 9035 -138 9135 -100
rect 9035 -172 9051 -138
rect 9119 -172 9135 -138
rect 9035 -188 9135 -172
rect 9193 -138 9293 -100
rect 9193 -172 9209 -138
rect 9277 -172 9293 -138
rect 9193 -188 9293 -172
rect 9351 -138 9451 -100
rect 9351 -172 9367 -138
rect 9435 -172 9451 -138
rect 9351 -188 9451 -172
<< polycont >>
rect -9435 138 -9367 172
rect -9277 138 -9209 172
rect -9119 138 -9051 172
rect -8961 138 -8893 172
rect -8803 138 -8735 172
rect -8645 138 -8577 172
rect -8487 138 -8419 172
rect -8329 138 -8261 172
rect -8171 138 -8103 172
rect -8013 138 -7945 172
rect -7855 138 -7787 172
rect -7697 138 -7629 172
rect -7539 138 -7471 172
rect -7381 138 -7313 172
rect -7223 138 -7155 172
rect -7065 138 -6997 172
rect -6907 138 -6839 172
rect -6749 138 -6681 172
rect -6591 138 -6523 172
rect -6433 138 -6365 172
rect -6275 138 -6207 172
rect -6117 138 -6049 172
rect -5959 138 -5891 172
rect -5801 138 -5733 172
rect -5643 138 -5575 172
rect -5485 138 -5417 172
rect -5327 138 -5259 172
rect -5169 138 -5101 172
rect -5011 138 -4943 172
rect -4853 138 -4785 172
rect -4695 138 -4627 172
rect -4537 138 -4469 172
rect -4379 138 -4311 172
rect -4221 138 -4153 172
rect -4063 138 -3995 172
rect -3905 138 -3837 172
rect -3747 138 -3679 172
rect -3589 138 -3521 172
rect -3431 138 -3363 172
rect -3273 138 -3205 172
rect -3115 138 -3047 172
rect -2957 138 -2889 172
rect -2799 138 -2731 172
rect -2641 138 -2573 172
rect -2483 138 -2415 172
rect -2325 138 -2257 172
rect -2167 138 -2099 172
rect -2009 138 -1941 172
rect -1851 138 -1783 172
rect -1693 138 -1625 172
rect -1535 138 -1467 172
rect -1377 138 -1309 172
rect -1219 138 -1151 172
rect -1061 138 -993 172
rect -903 138 -835 172
rect -745 138 -677 172
rect -587 138 -519 172
rect -429 138 -361 172
rect -271 138 -203 172
rect -113 138 -45 172
rect 45 138 113 172
rect 203 138 271 172
rect 361 138 429 172
rect 519 138 587 172
rect 677 138 745 172
rect 835 138 903 172
rect 993 138 1061 172
rect 1151 138 1219 172
rect 1309 138 1377 172
rect 1467 138 1535 172
rect 1625 138 1693 172
rect 1783 138 1851 172
rect 1941 138 2009 172
rect 2099 138 2167 172
rect 2257 138 2325 172
rect 2415 138 2483 172
rect 2573 138 2641 172
rect 2731 138 2799 172
rect 2889 138 2957 172
rect 3047 138 3115 172
rect 3205 138 3273 172
rect 3363 138 3431 172
rect 3521 138 3589 172
rect 3679 138 3747 172
rect 3837 138 3905 172
rect 3995 138 4063 172
rect 4153 138 4221 172
rect 4311 138 4379 172
rect 4469 138 4537 172
rect 4627 138 4695 172
rect 4785 138 4853 172
rect 4943 138 5011 172
rect 5101 138 5169 172
rect 5259 138 5327 172
rect 5417 138 5485 172
rect 5575 138 5643 172
rect 5733 138 5801 172
rect 5891 138 5959 172
rect 6049 138 6117 172
rect 6207 138 6275 172
rect 6365 138 6433 172
rect 6523 138 6591 172
rect 6681 138 6749 172
rect 6839 138 6907 172
rect 6997 138 7065 172
rect 7155 138 7223 172
rect 7313 138 7381 172
rect 7471 138 7539 172
rect 7629 138 7697 172
rect 7787 138 7855 172
rect 7945 138 8013 172
rect 8103 138 8171 172
rect 8261 138 8329 172
rect 8419 138 8487 172
rect 8577 138 8645 172
rect 8735 138 8803 172
rect 8893 138 8961 172
rect 9051 138 9119 172
rect 9209 138 9277 172
rect 9367 138 9435 172
rect -9435 -172 -9367 -138
rect -9277 -172 -9209 -138
rect -9119 -172 -9051 -138
rect -8961 -172 -8893 -138
rect -8803 -172 -8735 -138
rect -8645 -172 -8577 -138
rect -8487 -172 -8419 -138
rect -8329 -172 -8261 -138
rect -8171 -172 -8103 -138
rect -8013 -172 -7945 -138
rect -7855 -172 -7787 -138
rect -7697 -172 -7629 -138
rect -7539 -172 -7471 -138
rect -7381 -172 -7313 -138
rect -7223 -172 -7155 -138
rect -7065 -172 -6997 -138
rect -6907 -172 -6839 -138
rect -6749 -172 -6681 -138
rect -6591 -172 -6523 -138
rect -6433 -172 -6365 -138
rect -6275 -172 -6207 -138
rect -6117 -172 -6049 -138
rect -5959 -172 -5891 -138
rect -5801 -172 -5733 -138
rect -5643 -172 -5575 -138
rect -5485 -172 -5417 -138
rect -5327 -172 -5259 -138
rect -5169 -172 -5101 -138
rect -5011 -172 -4943 -138
rect -4853 -172 -4785 -138
rect -4695 -172 -4627 -138
rect -4537 -172 -4469 -138
rect -4379 -172 -4311 -138
rect -4221 -172 -4153 -138
rect -4063 -172 -3995 -138
rect -3905 -172 -3837 -138
rect -3747 -172 -3679 -138
rect -3589 -172 -3521 -138
rect -3431 -172 -3363 -138
rect -3273 -172 -3205 -138
rect -3115 -172 -3047 -138
rect -2957 -172 -2889 -138
rect -2799 -172 -2731 -138
rect -2641 -172 -2573 -138
rect -2483 -172 -2415 -138
rect -2325 -172 -2257 -138
rect -2167 -172 -2099 -138
rect -2009 -172 -1941 -138
rect -1851 -172 -1783 -138
rect -1693 -172 -1625 -138
rect -1535 -172 -1467 -138
rect -1377 -172 -1309 -138
rect -1219 -172 -1151 -138
rect -1061 -172 -993 -138
rect -903 -172 -835 -138
rect -745 -172 -677 -138
rect -587 -172 -519 -138
rect -429 -172 -361 -138
rect -271 -172 -203 -138
rect -113 -172 -45 -138
rect 45 -172 113 -138
rect 203 -172 271 -138
rect 361 -172 429 -138
rect 519 -172 587 -138
rect 677 -172 745 -138
rect 835 -172 903 -138
rect 993 -172 1061 -138
rect 1151 -172 1219 -138
rect 1309 -172 1377 -138
rect 1467 -172 1535 -138
rect 1625 -172 1693 -138
rect 1783 -172 1851 -138
rect 1941 -172 2009 -138
rect 2099 -172 2167 -138
rect 2257 -172 2325 -138
rect 2415 -172 2483 -138
rect 2573 -172 2641 -138
rect 2731 -172 2799 -138
rect 2889 -172 2957 -138
rect 3047 -172 3115 -138
rect 3205 -172 3273 -138
rect 3363 -172 3431 -138
rect 3521 -172 3589 -138
rect 3679 -172 3747 -138
rect 3837 -172 3905 -138
rect 3995 -172 4063 -138
rect 4153 -172 4221 -138
rect 4311 -172 4379 -138
rect 4469 -172 4537 -138
rect 4627 -172 4695 -138
rect 4785 -172 4853 -138
rect 4943 -172 5011 -138
rect 5101 -172 5169 -138
rect 5259 -172 5327 -138
rect 5417 -172 5485 -138
rect 5575 -172 5643 -138
rect 5733 -172 5801 -138
rect 5891 -172 5959 -138
rect 6049 -172 6117 -138
rect 6207 -172 6275 -138
rect 6365 -172 6433 -138
rect 6523 -172 6591 -138
rect 6681 -172 6749 -138
rect 6839 -172 6907 -138
rect 6997 -172 7065 -138
rect 7155 -172 7223 -138
rect 7313 -172 7381 -138
rect 7471 -172 7539 -138
rect 7629 -172 7697 -138
rect 7787 -172 7855 -138
rect 7945 -172 8013 -138
rect 8103 -172 8171 -138
rect 8261 -172 8329 -138
rect 8419 -172 8487 -138
rect 8577 -172 8645 -138
rect 8735 -172 8803 -138
rect 8893 -172 8961 -138
rect 9051 -172 9119 -138
rect 9209 -172 9277 -138
rect 9367 -172 9435 -138
<< locali >>
rect -9631 276 -9535 310
rect 9535 276 9631 310
rect -9631 214 -9597 276
rect 9597 214 9631 276
rect -9451 138 -9435 172
rect -9367 138 -9351 172
rect -9293 138 -9277 172
rect -9209 138 -9193 172
rect -9135 138 -9119 172
rect -9051 138 -9035 172
rect -8977 138 -8961 172
rect -8893 138 -8877 172
rect -8819 138 -8803 172
rect -8735 138 -8719 172
rect -8661 138 -8645 172
rect -8577 138 -8561 172
rect -8503 138 -8487 172
rect -8419 138 -8403 172
rect -8345 138 -8329 172
rect -8261 138 -8245 172
rect -8187 138 -8171 172
rect -8103 138 -8087 172
rect -8029 138 -8013 172
rect -7945 138 -7929 172
rect -7871 138 -7855 172
rect -7787 138 -7771 172
rect -7713 138 -7697 172
rect -7629 138 -7613 172
rect -7555 138 -7539 172
rect -7471 138 -7455 172
rect -7397 138 -7381 172
rect -7313 138 -7297 172
rect -7239 138 -7223 172
rect -7155 138 -7139 172
rect -7081 138 -7065 172
rect -6997 138 -6981 172
rect -6923 138 -6907 172
rect -6839 138 -6823 172
rect -6765 138 -6749 172
rect -6681 138 -6665 172
rect -6607 138 -6591 172
rect -6523 138 -6507 172
rect -6449 138 -6433 172
rect -6365 138 -6349 172
rect -6291 138 -6275 172
rect -6207 138 -6191 172
rect -6133 138 -6117 172
rect -6049 138 -6033 172
rect -5975 138 -5959 172
rect -5891 138 -5875 172
rect -5817 138 -5801 172
rect -5733 138 -5717 172
rect -5659 138 -5643 172
rect -5575 138 -5559 172
rect -5501 138 -5485 172
rect -5417 138 -5401 172
rect -5343 138 -5327 172
rect -5259 138 -5243 172
rect -5185 138 -5169 172
rect -5101 138 -5085 172
rect -5027 138 -5011 172
rect -4943 138 -4927 172
rect -4869 138 -4853 172
rect -4785 138 -4769 172
rect -4711 138 -4695 172
rect -4627 138 -4611 172
rect -4553 138 -4537 172
rect -4469 138 -4453 172
rect -4395 138 -4379 172
rect -4311 138 -4295 172
rect -4237 138 -4221 172
rect -4153 138 -4137 172
rect -4079 138 -4063 172
rect -3995 138 -3979 172
rect -3921 138 -3905 172
rect -3837 138 -3821 172
rect -3763 138 -3747 172
rect -3679 138 -3663 172
rect -3605 138 -3589 172
rect -3521 138 -3505 172
rect -3447 138 -3431 172
rect -3363 138 -3347 172
rect -3289 138 -3273 172
rect -3205 138 -3189 172
rect -3131 138 -3115 172
rect -3047 138 -3031 172
rect -2973 138 -2957 172
rect -2889 138 -2873 172
rect -2815 138 -2799 172
rect -2731 138 -2715 172
rect -2657 138 -2641 172
rect -2573 138 -2557 172
rect -2499 138 -2483 172
rect -2415 138 -2399 172
rect -2341 138 -2325 172
rect -2257 138 -2241 172
rect -2183 138 -2167 172
rect -2099 138 -2083 172
rect -2025 138 -2009 172
rect -1941 138 -1925 172
rect -1867 138 -1851 172
rect -1783 138 -1767 172
rect -1709 138 -1693 172
rect -1625 138 -1609 172
rect -1551 138 -1535 172
rect -1467 138 -1451 172
rect -1393 138 -1377 172
rect -1309 138 -1293 172
rect -1235 138 -1219 172
rect -1151 138 -1135 172
rect -1077 138 -1061 172
rect -993 138 -977 172
rect -919 138 -903 172
rect -835 138 -819 172
rect -761 138 -745 172
rect -677 138 -661 172
rect -603 138 -587 172
rect -519 138 -503 172
rect -445 138 -429 172
rect -361 138 -345 172
rect -287 138 -271 172
rect -203 138 -187 172
rect -129 138 -113 172
rect -45 138 -29 172
rect 29 138 45 172
rect 113 138 129 172
rect 187 138 203 172
rect 271 138 287 172
rect 345 138 361 172
rect 429 138 445 172
rect 503 138 519 172
rect 587 138 603 172
rect 661 138 677 172
rect 745 138 761 172
rect 819 138 835 172
rect 903 138 919 172
rect 977 138 993 172
rect 1061 138 1077 172
rect 1135 138 1151 172
rect 1219 138 1235 172
rect 1293 138 1309 172
rect 1377 138 1393 172
rect 1451 138 1467 172
rect 1535 138 1551 172
rect 1609 138 1625 172
rect 1693 138 1709 172
rect 1767 138 1783 172
rect 1851 138 1867 172
rect 1925 138 1941 172
rect 2009 138 2025 172
rect 2083 138 2099 172
rect 2167 138 2183 172
rect 2241 138 2257 172
rect 2325 138 2341 172
rect 2399 138 2415 172
rect 2483 138 2499 172
rect 2557 138 2573 172
rect 2641 138 2657 172
rect 2715 138 2731 172
rect 2799 138 2815 172
rect 2873 138 2889 172
rect 2957 138 2973 172
rect 3031 138 3047 172
rect 3115 138 3131 172
rect 3189 138 3205 172
rect 3273 138 3289 172
rect 3347 138 3363 172
rect 3431 138 3447 172
rect 3505 138 3521 172
rect 3589 138 3605 172
rect 3663 138 3679 172
rect 3747 138 3763 172
rect 3821 138 3837 172
rect 3905 138 3921 172
rect 3979 138 3995 172
rect 4063 138 4079 172
rect 4137 138 4153 172
rect 4221 138 4237 172
rect 4295 138 4311 172
rect 4379 138 4395 172
rect 4453 138 4469 172
rect 4537 138 4553 172
rect 4611 138 4627 172
rect 4695 138 4711 172
rect 4769 138 4785 172
rect 4853 138 4869 172
rect 4927 138 4943 172
rect 5011 138 5027 172
rect 5085 138 5101 172
rect 5169 138 5185 172
rect 5243 138 5259 172
rect 5327 138 5343 172
rect 5401 138 5417 172
rect 5485 138 5501 172
rect 5559 138 5575 172
rect 5643 138 5659 172
rect 5717 138 5733 172
rect 5801 138 5817 172
rect 5875 138 5891 172
rect 5959 138 5975 172
rect 6033 138 6049 172
rect 6117 138 6133 172
rect 6191 138 6207 172
rect 6275 138 6291 172
rect 6349 138 6365 172
rect 6433 138 6449 172
rect 6507 138 6523 172
rect 6591 138 6607 172
rect 6665 138 6681 172
rect 6749 138 6765 172
rect 6823 138 6839 172
rect 6907 138 6923 172
rect 6981 138 6997 172
rect 7065 138 7081 172
rect 7139 138 7155 172
rect 7223 138 7239 172
rect 7297 138 7313 172
rect 7381 138 7397 172
rect 7455 138 7471 172
rect 7539 138 7555 172
rect 7613 138 7629 172
rect 7697 138 7713 172
rect 7771 138 7787 172
rect 7855 138 7871 172
rect 7929 138 7945 172
rect 8013 138 8029 172
rect 8087 138 8103 172
rect 8171 138 8187 172
rect 8245 138 8261 172
rect 8329 138 8345 172
rect 8403 138 8419 172
rect 8487 138 8503 172
rect 8561 138 8577 172
rect 8645 138 8661 172
rect 8719 138 8735 172
rect 8803 138 8819 172
rect 8877 138 8893 172
rect 8961 138 8977 172
rect 9035 138 9051 172
rect 9119 138 9135 172
rect 9193 138 9209 172
rect 9277 138 9293 172
rect 9351 138 9367 172
rect 9435 138 9451 172
rect -9497 88 -9463 104
rect -9497 -104 -9463 -88
rect -9339 88 -9305 104
rect -9339 -104 -9305 -88
rect -9181 88 -9147 104
rect -9181 -104 -9147 -88
rect -9023 88 -8989 104
rect -9023 -104 -8989 -88
rect -8865 88 -8831 104
rect -8865 -104 -8831 -88
rect -8707 88 -8673 104
rect -8707 -104 -8673 -88
rect -8549 88 -8515 104
rect -8549 -104 -8515 -88
rect -8391 88 -8357 104
rect -8391 -104 -8357 -88
rect -8233 88 -8199 104
rect -8233 -104 -8199 -88
rect -8075 88 -8041 104
rect -8075 -104 -8041 -88
rect -7917 88 -7883 104
rect -7917 -104 -7883 -88
rect -7759 88 -7725 104
rect -7759 -104 -7725 -88
rect -7601 88 -7567 104
rect -7601 -104 -7567 -88
rect -7443 88 -7409 104
rect -7443 -104 -7409 -88
rect -7285 88 -7251 104
rect -7285 -104 -7251 -88
rect -7127 88 -7093 104
rect -7127 -104 -7093 -88
rect -6969 88 -6935 104
rect -6969 -104 -6935 -88
rect -6811 88 -6777 104
rect -6811 -104 -6777 -88
rect -6653 88 -6619 104
rect -6653 -104 -6619 -88
rect -6495 88 -6461 104
rect -6495 -104 -6461 -88
rect -6337 88 -6303 104
rect -6337 -104 -6303 -88
rect -6179 88 -6145 104
rect -6179 -104 -6145 -88
rect -6021 88 -5987 104
rect -6021 -104 -5987 -88
rect -5863 88 -5829 104
rect -5863 -104 -5829 -88
rect -5705 88 -5671 104
rect -5705 -104 -5671 -88
rect -5547 88 -5513 104
rect -5547 -104 -5513 -88
rect -5389 88 -5355 104
rect -5389 -104 -5355 -88
rect -5231 88 -5197 104
rect -5231 -104 -5197 -88
rect -5073 88 -5039 104
rect -5073 -104 -5039 -88
rect -4915 88 -4881 104
rect -4915 -104 -4881 -88
rect -4757 88 -4723 104
rect -4757 -104 -4723 -88
rect -4599 88 -4565 104
rect -4599 -104 -4565 -88
rect -4441 88 -4407 104
rect -4441 -104 -4407 -88
rect -4283 88 -4249 104
rect -4283 -104 -4249 -88
rect -4125 88 -4091 104
rect -4125 -104 -4091 -88
rect -3967 88 -3933 104
rect -3967 -104 -3933 -88
rect -3809 88 -3775 104
rect -3809 -104 -3775 -88
rect -3651 88 -3617 104
rect -3651 -104 -3617 -88
rect -3493 88 -3459 104
rect -3493 -104 -3459 -88
rect -3335 88 -3301 104
rect -3335 -104 -3301 -88
rect -3177 88 -3143 104
rect -3177 -104 -3143 -88
rect -3019 88 -2985 104
rect -3019 -104 -2985 -88
rect -2861 88 -2827 104
rect -2861 -104 -2827 -88
rect -2703 88 -2669 104
rect -2703 -104 -2669 -88
rect -2545 88 -2511 104
rect -2545 -104 -2511 -88
rect -2387 88 -2353 104
rect -2387 -104 -2353 -88
rect -2229 88 -2195 104
rect -2229 -104 -2195 -88
rect -2071 88 -2037 104
rect -2071 -104 -2037 -88
rect -1913 88 -1879 104
rect -1913 -104 -1879 -88
rect -1755 88 -1721 104
rect -1755 -104 -1721 -88
rect -1597 88 -1563 104
rect -1597 -104 -1563 -88
rect -1439 88 -1405 104
rect -1439 -104 -1405 -88
rect -1281 88 -1247 104
rect -1281 -104 -1247 -88
rect -1123 88 -1089 104
rect -1123 -104 -1089 -88
rect -965 88 -931 104
rect -965 -104 -931 -88
rect -807 88 -773 104
rect -807 -104 -773 -88
rect -649 88 -615 104
rect -649 -104 -615 -88
rect -491 88 -457 104
rect -491 -104 -457 -88
rect -333 88 -299 104
rect -333 -104 -299 -88
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect 299 88 333 104
rect 299 -104 333 -88
rect 457 88 491 104
rect 457 -104 491 -88
rect 615 88 649 104
rect 615 -104 649 -88
rect 773 88 807 104
rect 773 -104 807 -88
rect 931 88 965 104
rect 931 -104 965 -88
rect 1089 88 1123 104
rect 1089 -104 1123 -88
rect 1247 88 1281 104
rect 1247 -104 1281 -88
rect 1405 88 1439 104
rect 1405 -104 1439 -88
rect 1563 88 1597 104
rect 1563 -104 1597 -88
rect 1721 88 1755 104
rect 1721 -104 1755 -88
rect 1879 88 1913 104
rect 1879 -104 1913 -88
rect 2037 88 2071 104
rect 2037 -104 2071 -88
rect 2195 88 2229 104
rect 2195 -104 2229 -88
rect 2353 88 2387 104
rect 2353 -104 2387 -88
rect 2511 88 2545 104
rect 2511 -104 2545 -88
rect 2669 88 2703 104
rect 2669 -104 2703 -88
rect 2827 88 2861 104
rect 2827 -104 2861 -88
rect 2985 88 3019 104
rect 2985 -104 3019 -88
rect 3143 88 3177 104
rect 3143 -104 3177 -88
rect 3301 88 3335 104
rect 3301 -104 3335 -88
rect 3459 88 3493 104
rect 3459 -104 3493 -88
rect 3617 88 3651 104
rect 3617 -104 3651 -88
rect 3775 88 3809 104
rect 3775 -104 3809 -88
rect 3933 88 3967 104
rect 3933 -104 3967 -88
rect 4091 88 4125 104
rect 4091 -104 4125 -88
rect 4249 88 4283 104
rect 4249 -104 4283 -88
rect 4407 88 4441 104
rect 4407 -104 4441 -88
rect 4565 88 4599 104
rect 4565 -104 4599 -88
rect 4723 88 4757 104
rect 4723 -104 4757 -88
rect 4881 88 4915 104
rect 4881 -104 4915 -88
rect 5039 88 5073 104
rect 5039 -104 5073 -88
rect 5197 88 5231 104
rect 5197 -104 5231 -88
rect 5355 88 5389 104
rect 5355 -104 5389 -88
rect 5513 88 5547 104
rect 5513 -104 5547 -88
rect 5671 88 5705 104
rect 5671 -104 5705 -88
rect 5829 88 5863 104
rect 5829 -104 5863 -88
rect 5987 88 6021 104
rect 5987 -104 6021 -88
rect 6145 88 6179 104
rect 6145 -104 6179 -88
rect 6303 88 6337 104
rect 6303 -104 6337 -88
rect 6461 88 6495 104
rect 6461 -104 6495 -88
rect 6619 88 6653 104
rect 6619 -104 6653 -88
rect 6777 88 6811 104
rect 6777 -104 6811 -88
rect 6935 88 6969 104
rect 6935 -104 6969 -88
rect 7093 88 7127 104
rect 7093 -104 7127 -88
rect 7251 88 7285 104
rect 7251 -104 7285 -88
rect 7409 88 7443 104
rect 7409 -104 7443 -88
rect 7567 88 7601 104
rect 7567 -104 7601 -88
rect 7725 88 7759 104
rect 7725 -104 7759 -88
rect 7883 88 7917 104
rect 7883 -104 7917 -88
rect 8041 88 8075 104
rect 8041 -104 8075 -88
rect 8199 88 8233 104
rect 8199 -104 8233 -88
rect 8357 88 8391 104
rect 8357 -104 8391 -88
rect 8515 88 8549 104
rect 8515 -104 8549 -88
rect 8673 88 8707 104
rect 8673 -104 8707 -88
rect 8831 88 8865 104
rect 8831 -104 8865 -88
rect 8989 88 9023 104
rect 8989 -104 9023 -88
rect 9147 88 9181 104
rect 9147 -104 9181 -88
rect 9305 88 9339 104
rect 9305 -104 9339 -88
rect 9463 88 9497 104
rect 9463 -104 9497 -88
rect -9451 -172 -9435 -138
rect -9367 -172 -9351 -138
rect -9293 -172 -9277 -138
rect -9209 -172 -9193 -138
rect -9135 -172 -9119 -138
rect -9051 -172 -9035 -138
rect -8977 -172 -8961 -138
rect -8893 -172 -8877 -138
rect -8819 -172 -8803 -138
rect -8735 -172 -8719 -138
rect -8661 -172 -8645 -138
rect -8577 -172 -8561 -138
rect -8503 -172 -8487 -138
rect -8419 -172 -8403 -138
rect -8345 -172 -8329 -138
rect -8261 -172 -8245 -138
rect -8187 -172 -8171 -138
rect -8103 -172 -8087 -138
rect -8029 -172 -8013 -138
rect -7945 -172 -7929 -138
rect -7871 -172 -7855 -138
rect -7787 -172 -7771 -138
rect -7713 -172 -7697 -138
rect -7629 -172 -7613 -138
rect -7555 -172 -7539 -138
rect -7471 -172 -7455 -138
rect -7397 -172 -7381 -138
rect -7313 -172 -7297 -138
rect -7239 -172 -7223 -138
rect -7155 -172 -7139 -138
rect -7081 -172 -7065 -138
rect -6997 -172 -6981 -138
rect -6923 -172 -6907 -138
rect -6839 -172 -6823 -138
rect -6765 -172 -6749 -138
rect -6681 -172 -6665 -138
rect -6607 -172 -6591 -138
rect -6523 -172 -6507 -138
rect -6449 -172 -6433 -138
rect -6365 -172 -6349 -138
rect -6291 -172 -6275 -138
rect -6207 -172 -6191 -138
rect -6133 -172 -6117 -138
rect -6049 -172 -6033 -138
rect -5975 -172 -5959 -138
rect -5891 -172 -5875 -138
rect -5817 -172 -5801 -138
rect -5733 -172 -5717 -138
rect -5659 -172 -5643 -138
rect -5575 -172 -5559 -138
rect -5501 -172 -5485 -138
rect -5417 -172 -5401 -138
rect -5343 -172 -5327 -138
rect -5259 -172 -5243 -138
rect -5185 -172 -5169 -138
rect -5101 -172 -5085 -138
rect -5027 -172 -5011 -138
rect -4943 -172 -4927 -138
rect -4869 -172 -4853 -138
rect -4785 -172 -4769 -138
rect -4711 -172 -4695 -138
rect -4627 -172 -4611 -138
rect -4553 -172 -4537 -138
rect -4469 -172 -4453 -138
rect -4395 -172 -4379 -138
rect -4311 -172 -4295 -138
rect -4237 -172 -4221 -138
rect -4153 -172 -4137 -138
rect -4079 -172 -4063 -138
rect -3995 -172 -3979 -138
rect -3921 -172 -3905 -138
rect -3837 -172 -3821 -138
rect -3763 -172 -3747 -138
rect -3679 -172 -3663 -138
rect -3605 -172 -3589 -138
rect -3521 -172 -3505 -138
rect -3447 -172 -3431 -138
rect -3363 -172 -3347 -138
rect -3289 -172 -3273 -138
rect -3205 -172 -3189 -138
rect -3131 -172 -3115 -138
rect -3047 -172 -3031 -138
rect -2973 -172 -2957 -138
rect -2889 -172 -2873 -138
rect -2815 -172 -2799 -138
rect -2731 -172 -2715 -138
rect -2657 -172 -2641 -138
rect -2573 -172 -2557 -138
rect -2499 -172 -2483 -138
rect -2415 -172 -2399 -138
rect -2341 -172 -2325 -138
rect -2257 -172 -2241 -138
rect -2183 -172 -2167 -138
rect -2099 -172 -2083 -138
rect -2025 -172 -2009 -138
rect -1941 -172 -1925 -138
rect -1867 -172 -1851 -138
rect -1783 -172 -1767 -138
rect -1709 -172 -1693 -138
rect -1625 -172 -1609 -138
rect -1551 -172 -1535 -138
rect -1467 -172 -1451 -138
rect -1393 -172 -1377 -138
rect -1309 -172 -1293 -138
rect -1235 -172 -1219 -138
rect -1151 -172 -1135 -138
rect -1077 -172 -1061 -138
rect -993 -172 -977 -138
rect -919 -172 -903 -138
rect -835 -172 -819 -138
rect -761 -172 -745 -138
rect -677 -172 -661 -138
rect -603 -172 -587 -138
rect -519 -172 -503 -138
rect -445 -172 -429 -138
rect -361 -172 -345 -138
rect -287 -172 -271 -138
rect -203 -172 -187 -138
rect -129 -172 -113 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 113 -172 129 -138
rect 187 -172 203 -138
rect 271 -172 287 -138
rect 345 -172 361 -138
rect 429 -172 445 -138
rect 503 -172 519 -138
rect 587 -172 603 -138
rect 661 -172 677 -138
rect 745 -172 761 -138
rect 819 -172 835 -138
rect 903 -172 919 -138
rect 977 -172 993 -138
rect 1061 -172 1077 -138
rect 1135 -172 1151 -138
rect 1219 -172 1235 -138
rect 1293 -172 1309 -138
rect 1377 -172 1393 -138
rect 1451 -172 1467 -138
rect 1535 -172 1551 -138
rect 1609 -172 1625 -138
rect 1693 -172 1709 -138
rect 1767 -172 1783 -138
rect 1851 -172 1867 -138
rect 1925 -172 1941 -138
rect 2009 -172 2025 -138
rect 2083 -172 2099 -138
rect 2167 -172 2183 -138
rect 2241 -172 2257 -138
rect 2325 -172 2341 -138
rect 2399 -172 2415 -138
rect 2483 -172 2499 -138
rect 2557 -172 2573 -138
rect 2641 -172 2657 -138
rect 2715 -172 2731 -138
rect 2799 -172 2815 -138
rect 2873 -172 2889 -138
rect 2957 -172 2973 -138
rect 3031 -172 3047 -138
rect 3115 -172 3131 -138
rect 3189 -172 3205 -138
rect 3273 -172 3289 -138
rect 3347 -172 3363 -138
rect 3431 -172 3447 -138
rect 3505 -172 3521 -138
rect 3589 -172 3605 -138
rect 3663 -172 3679 -138
rect 3747 -172 3763 -138
rect 3821 -172 3837 -138
rect 3905 -172 3921 -138
rect 3979 -172 3995 -138
rect 4063 -172 4079 -138
rect 4137 -172 4153 -138
rect 4221 -172 4237 -138
rect 4295 -172 4311 -138
rect 4379 -172 4395 -138
rect 4453 -172 4469 -138
rect 4537 -172 4553 -138
rect 4611 -172 4627 -138
rect 4695 -172 4711 -138
rect 4769 -172 4785 -138
rect 4853 -172 4869 -138
rect 4927 -172 4943 -138
rect 5011 -172 5027 -138
rect 5085 -172 5101 -138
rect 5169 -172 5185 -138
rect 5243 -172 5259 -138
rect 5327 -172 5343 -138
rect 5401 -172 5417 -138
rect 5485 -172 5501 -138
rect 5559 -172 5575 -138
rect 5643 -172 5659 -138
rect 5717 -172 5733 -138
rect 5801 -172 5817 -138
rect 5875 -172 5891 -138
rect 5959 -172 5975 -138
rect 6033 -172 6049 -138
rect 6117 -172 6133 -138
rect 6191 -172 6207 -138
rect 6275 -172 6291 -138
rect 6349 -172 6365 -138
rect 6433 -172 6449 -138
rect 6507 -172 6523 -138
rect 6591 -172 6607 -138
rect 6665 -172 6681 -138
rect 6749 -172 6765 -138
rect 6823 -172 6839 -138
rect 6907 -172 6923 -138
rect 6981 -172 6997 -138
rect 7065 -172 7081 -138
rect 7139 -172 7155 -138
rect 7223 -172 7239 -138
rect 7297 -172 7313 -138
rect 7381 -172 7397 -138
rect 7455 -172 7471 -138
rect 7539 -172 7555 -138
rect 7613 -172 7629 -138
rect 7697 -172 7713 -138
rect 7771 -172 7787 -138
rect 7855 -172 7871 -138
rect 7929 -172 7945 -138
rect 8013 -172 8029 -138
rect 8087 -172 8103 -138
rect 8171 -172 8187 -138
rect 8245 -172 8261 -138
rect 8329 -172 8345 -138
rect 8403 -172 8419 -138
rect 8487 -172 8503 -138
rect 8561 -172 8577 -138
rect 8645 -172 8661 -138
rect 8719 -172 8735 -138
rect 8803 -172 8819 -138
rect 8877 -172 8893 -138
rect 8961 -172 8977 -138
rect 9035 -172 9051 -138
rect 9119 -172 9135 -138
rect 9193 -172 9209 -138
rect 9277 -172 9293 -138
rect 9351 -172 9367 -138
rect 9435 -172 9451 -138
rect -9631 -276 -9597 -214
rect 9597 -276 9631 -214
rect -9631 -310 -9535 -276
rect 9535 -310 9631 -276
<< viali >>
rect -9435 138 -9367 172
rect -9277 138 -9209 172
rect -9119 138 -9051 172
rect -8961 138 -8893 172
rect -8803 138 -8735 172
rect -8645 138 -8577 172
rect -8487 138 -8419 172
rect -8329 138 -8261 172
rect -8171 138 -8103 172
rect -8013 138 -7945 172
rect -7855 138 -7787 172
rect -7697 138 -7629 172
rect -7539 138 -7471 172
rect -7381 138 -7313 172
rect -7223 138 -7155 172
rect -7065 138 -6997 172
rect -6907 138 -6839 172
rect -6749 138 -6681 172
rect -6591 138 -6523 172
rect -6433 138 -6365 172
rect -6275 138 -6207 172
rect -6117 138 -6049 172
rect -5959 138 -5891 172
rect -5801 138 -5733 172
rect -5643 138 -5575 172
rect -5485 138 -5417 172
rect -5327 138 -5259 172
rect -5169 138 -5101 172
rect -5011 138 -4943 172
rect -4853 138 -4785 172
rect -4695 138 -4627 172
rect -4537 138 -4469 172
rect -4379 138 -4311 172
rect -4221 138 -4153 172
rect -4063 138 -3995 172
rect -3905 138 -3837 172
rect -3747 138 -3679 172
rect -3589 138 -3521 172
rect -3431 138 -3363 172
rect -3273 138 -3205 172
rect -3115 138 -3047 172
rect -2957 138 -2889 172
rect -2799 138 -2731 172
rect -2641 138 -2573 172
rect -2483 138 -2415 172
rect -2325 138 -2257 172
rect -2167 138 -2099 172
rect -2009 138 -1941 172
rect -1851 138 -1783 172
rect -1693 138 -1625 172
rect -1535 138 -1467 172
rect -1377 138 -1309 172
rect -1219 138 -1151 172
rect -1061 138 -993 172
rect -903 138 -835 172
rect -745 138 -677 172
rect -587 138 -519 172
rect -429 138 -361 172
rect -271 138 -203 172
rect -113 138 -45 172
rect 45 138 113 172
rect 203 138 271 172
rect 361 138 429 172
rect 519 138 587 172
rect 677 138 745 172
rect 835 138 903 172
rect 993 138 1061 172
rect 1151 138 1219 172
rect 1309 138 1377 172
rect 1467 138 1535 172
rect 1625 138 1693 172
rect 1783 138 1851 172
rect 1941 138 2009 172
rect 2099 138 2167 172
rect 2257 138 2325 172
rect 2415 138 2483 172
rect 2573 138 2641 172
rect 2731 138 2799 172
rect 2889 138 2957 172
rect 3047 138 3115 172
rect 3205 138 3273 172
rect 3363 138 3431 172
rect 3521 138 3589 172
rect 3679 138 3747 172
rect 3837 138 3905 172
rect 3995 138 4063 172
rect 4153 138 4221 172
rect 4311 138 4379 172
rect 4469 138 4537 172
rect 4627 138 4695 172
rect 4785 138 4853 172
rect 4943 138 5011 172
rect 5101 138 5169 172
rect 5259 138 5327 172
rect 5417 138 5485 172
rect 5575 138 5643 172
rect 5733 138 5801 172
rect 5891 138 5959 172
rect 6049 138 6117 172
rect 6207 138 6275 172
rect 6365 138 6433 172
rect 6523 138 6591 172
rect 6681 138 6749 172
rect 6839 138 6907 172
rect 6997 138 7065 172
rect 7155 138 7223 172
rect 7313 138 7381 172
rect 7471 138 7539 172
rect 7629 138 7697 172
rect 7787 138 7855 172
rect 7945 138 8013 172
rect 8103 138 8171 172
rect 8261 138 8329 172
rect 8419 138 8487 172
rect 8577 138 8645 172
rect 8735 138 8803 172
rect 8893 138 8961 172
rect 9051 138 9119 172
rect 9209 138 9277 172
rect 9367 138 9435 172
rect -9497 -88 -9463 88
rect -9339 -88 -9305 88
rect -9181 -88 -9147 88
rect -9023 -88 -8989 88
rect -8865 -88 -8831 88
rect -8707 -88 -8673 88
rect -8549 -88 -8515 88
rect -8391 -88 -8357 88
rect -8233 -88 -8199 88
rect -8075 -88 -8041 88
rect -7917 -88 -7883 88
rect -7759 -88 -7725 88
rect -7601 -88 -7567 88
rect -7443 -88 -7409 88
rect -7285 -88 -7251 88
rect -7127 -88 -7093 88
rect -6969 -88 -6935 88
rect -6811 -88 -6777 88
rect -6653 -88 -6619 88
rect -6495 -88 -6461 88
rect -6337 -88 -6303 88
rect -6179 -88 -6145 88
rect -6021 -88 -5987 88
rect -5863 -88 -5829 88
rect -5705 -88 -5671 88
rect -5547 -88 -5513 88
rect -5389 -88 -5355 88
rect -5231 -88 -5197 88
rect -5073 -88 -5039 88
rect -4915 -88 -4881 88
rect -4757 -88 -4723 88
rect -4599 -88 -4565 88
rect -4441 -88 -4407 88
rect -4283 -88 -4249 88
rect -4125 -88 -4091 88
rect -3967 -88 -3933 88
rect -3809 -88 -3775 88
rect -3651 -88 -3617 88
rect -3493 -88 -3459 88
rect -3335 -88 -3301 88
rect -3177 -88 -3143 88
rect -3019 -88 -2985 88
rect -2861 -88 -2827 88
rect -2703 -88 -2669 88
rect -2545 -88 -2511 88
rect -2387 -88 -2353 88
rect -2229 -88 -2195 88
rect -2071 -88 -2037 88
rect -1913 -88 -1879 88
rect -1755 -88 -1721 88
rect -1597 -88 -1563 88
rect -1439 -88 -1405 88
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
rect 1405 -88 1439 88
rect 1563 -88 1597 88
rect 1721 -88 1755 88
rect 1879 -88 1913 88
rect 2037 -88 2071 88
rect 2195 -88 2229 88
rect 2353 -88 2387 88
rect 2511 -88 2545 88
rect 2669 -88 2703 88
rect 2827 -88 2861 88
rect 2985 -88 3019 88
rect 3143 -88 3177 88
rect 3301 -88 3335 88
rect 3459 -88 3493 88
rect 3617 -88 3651 88
rect 3775 -88 3809 88
rect 3933 -88 3967 88
rect 4091 -88 4125 88
rect 4249 -88 4283 88
rect 4407 -88 4441 88
rect 4565 -88 4599 88
rect 4723 -88 4757 88
rect 4881 -88 4915 88
rect 5039 -88 5073 88
rect 5197 -88 5231 88
rect 5355 -88 5389 88
rect 5513 -88 5547 88
rect 5671 -88 5705 88
rect 5829 -88 5863 88
rect 5987 -88 6021 88
rect 6145 -88 6179 88
rect 6303 -88 6337 88
rect 6461 -88 6495 88
rect 6619 -88 6653 88
rect 6777 -88 6811 88
rect 6935 -88 6969 88
rect 7093 -88 7127 88
rect 7251 -88 7285 88
rect 7409 -88 7443 88
rect 7567 -88 7601 88
rect 7725 -88 7759 88
rect 7883 -88 7917 88
rect 8041 -88 8075 88
rect 8199 -88 8233 88
rect 8357 -88 8391 88
rect 8515 -88 8549 88
rect 8673 -88 8707 88
rect 8831 -88 8865 88
rect 8989 -88 9023 88
rect 9147 -88 9181 88
rect 9305 -88 9339 88
rect 9463 -88 9497 88
rect -9435 -172 -9367 -138
rect -9277 -172 -9209 -138
rect -9119 -172 -9051 -138
rect -8961 -172 -8893 -138
rect -8803 -172 -8735 -138
rect -8645 -172 -8577 -138
rect -8487 -172 -8419 -138
rect -8329 -172 -8261 -138
rect -8171 -172 -8103 -138
rect -8013 -172 -7945 -138
rect -7855 -172 -7787 -138
rect -7697 -172 -7629 -138
rect -7539 -172 -7471 -138
rect -7381 -172 -7313 -138
rect -7223 -172 -7155 -138
rect -7065 -172 -6997 -138
rect -6907 -172 -6839 -138
rect -6749 -172 -6681 -138
rect -6591 -172 -6523 -138
rect -6433 -172 -6365 -138
rect -6275 -172 -6207 -138
rect -6117 -172 -6049 -138
rect -5959 -172 -5891 -138
rect -5801 -172 -5733 -138
rect -5643 -172 -5575 -138
rect -5485 -172 -5417 -138
rect -5327 -172 -5259 -138
rect -5169 -172 -5101 -138
rect -5011 -172 -4943 -138
rect -4853 -172 -4785 -138
rect -4695 -172 -4627 -138
rect -4537 -172 -4469 -138
rect -4379 -172 -4311 -138
rect -4221 -172 -4153 -138
rect -4063 -172 -3995 -138
rect -3905 -172 -3837 -138
rect -3747 -172 -3679 -138
rect -3589 -172 -3521 -138
rect -3431 -172 -3363 -138
rect -3273 -172 -3205 -138
rect -3115 -172 -3047 -138
rect -2957 -172 -2889 -138
rect -2799 -172 -2731 -138
rect -2641 -172 -2573 -138
rect -2483 -172 -2415 -138
rect -2325 -172 -2257 -138
rect -2167 -172 -2099 -138
rect -2009 -172 -1941 -138
rect -1851 -172 -1783 -138
rect -1693 -172 -1625 -138
rect -1535 -172 -1467 -138
rect -1377 -172 -1309 -138
rect -1219 -172 -1151 -138
rect -1061 -172 -993 -138
rect -903 -172 -835 -138
rect -745 -172 -677 -138
rect -587 -172 -519 -138
rect -429 -172 -361 -138
rect -271 -172 -203 -138
rect -113 -172 -45 -138
rect 45 -172 113 -138
rect 203 -172 271 -138
rect 361 -172 429 -138
rect 519 -172 587 -138
rect 677 -172 745 -138
rect 835 -172 903 -138
rect 993 -172 1061 -138
rect 1151 -172 1219 -138
rect 1309 -172 1377 -138
rect 1467 -172 1535 -138
rect 1625 -172 1693 -138
rect 1783 -172 1851 -138
rect 1941 -172 2009 -138
rect 2099 -172 2167 -138
rect 2257 -172 2325 -138
rect 2415 -172 2483 -138
rect 2573 -172 2641 -138
rect 2731 -172 2799 -138
rect 2889 -172 2957 -138
rect 3047 -172 3115 -138
rect 3205 -172 3273 -138
rect 3363 -172 3431 -138
rect 3521 -172 3589 -138
rect 3679 -172 3747 -138
rect 3837 -172 3905 -138
rect 3995 -172 4063 -138
rect 4153 -172 4221 -138
rect 4311 -172 4379 -138
rect 4469 -172 4537 -138
rect 4627 -172 4695 -138
rect 4785 -172 4853 -138
rect 4943 -172 5011 -138
rect 5101 -172 5169 -138
rect 5259 -172 5327 -138
rect 5417 -172 5485 -138
rect 5575 -172 5643 -138
rect 5733 -172 5801 -138
rect 5891 -172 5959 -138
rect 6049 -172 6117 -138
rect 6207 -172 6275 -138
rect 6365 -172 6433 -138
rect 6523 -172 6591 -138
rect 6681 -172 6749 -138
rect 6839 -172 6907 -138
rect 6997 -172 7065 -138
rect 7155 -172 7223 -138
rect 7313 -172 7381 -138
rect 7471 -172 7539 -138
rect 7629 -172 7697 -138
rect 7787 -172 7855 -138
rect 7945 -172 8013 -138
rect 8103 -172 8171 -138
rect 8261 -172 8329 -138
rect 8419 -172 8487 -138
rect 8577 -172 8645 -138
rect 8735 -172 8803 -138
rect 8893 -172 8961 -138
rect 9051 -172 9119 -138
rect 9209 -172 9277 -138
rect 9367 -172 9435 -138
<< metal1 >>
rect -9447 172 -9355 178
rect -9447 138 -9435 172
rect -9367 138 -9355 172
rect -9447 132 -9355 138
rect -9289 172 -9197 178
rect -9289 138 -9277 172
rect -9209 138 -9197 172
rect -9289 132 -9197 138
rect -9131 172 -9039 178
rect -9131 138 -9119 172
rect -9051 138 -9039 172
rect -9131 132 -9039 138
rect -8973 172 -8881 178
rect -8973 138 -8961 172
rect -8893 138 -8881 172
rect -8973 132 -8881 138
rect -8815 172 -8723 178
rect -8815 138 -8803 172
rect -8735 138 -8723 172
rect -8815 132 -8723 138
rect -8657 172 -8565 178
rect -8657 138 -8645 172
rect -8577 138 -8565 172
rect -8657 132 -8565 138
rect -8499 172 -8407 178
rect -8499 138 -8487 172
rect -8419 138 -8407 172
rect -8499 132 -8407 138
rect -8341 172 -8249 178
rect -8341 138 -8329 172
rect -8261 138 -8249 172
rect -8341 132 -8249 138
rect -8183 172 -8091 178
rect -8183 138 -8171 172
rect -8103 138 -8091 172
rect -8183 132 -8091 138
rect -8025 172 -7933 178
rect -8025 138 -8013 172
rect -7945 138 -7933 172
rect -8025 132 -7933 138
rect -7867 172 -7775 178
rect -7867 138 -7855 172
rect -7787 138 -7775 172
rect -7867 132 -7775 138
rect -7709 172 -7617 178
rect -7709 138 -7697 172
rect -7629 138 -7617 172
rect -7709 132 -7617 138
rect -7551 172 -7459 178
rect -7551 138 -7539 172
rect -7471 138 -7459 172
rect -7551 132 -7459 138
rect -7393 172 -7301 178
rect -7393 138 -7381 172
rect -7313 138 -7301 172
rect -7393 132 -7301 138
rect -7235 172 -7143 178
rect -7235 138 -7223 172
rect -7155 138 -7143 172
rect -7235 132 -7143 138
rect -7077 172 -6985 178
rect -7077 138 -7065 172
rect -6997 138 -6985 172
rect -7077 132 -6985 138
rect -6919 172 -6827 178
rect -6919 138 -6907 172
rect -6839 138 -6827 172
rect -6919 132 -6827 138
rect -6761 172 -6669 178
rect -6761 138 -6749 172
rect -6681 138 -6669 172
rect -6761 132 -6669 138
rect -6603 172 -6511 178
rect -6603 138 -6591 172
rect -6523 138 -6511 172
rect -6603 132 -6511 138
rect -6445 172 -6353 178
rect -6445 138 -6433 172
rect -6365 138 -6353 172
rect -6445 132 -6353 138
rect -6287 172 -6195 178
rect -6287 138 -6275 172
rect -6207 138 -6195 172
rect -6287 132 -6195 138
rect -6129 172 -6037 178
rect -6129 138 -6117 172
rect -6049 138 -6037 172
rect -6129 132 -6037 138
rect -5971 172 -5879 178
rect -5971 138 -5959 172
rect -5891 138 -5879 172
rect -5971 132 -5879 138
rect -5813 172 -5721 178
rect -5813 138 -5801 172
rect -5733 138 -5721 172
rect -5813 132 -5721 138
rect -5655 172 -5563 178
rect -5655 138 -5643 172
rect -5575 138 -5563 172
rect -5655 132 -5563 138
rect -5497 172 -5405 178
rect -5497 138 -5485 172
rect -5417 138 -5405 172
rect -5497 132 -5405 138
rect -5339 172 -5247 178
rect -5339 138 -5327 172
rect -5259 138 -5247 172
rect -5339 132 -5247 138
rect -5181 172 -5089 178
rect -5181 138 -5169 172
rect -5101 138 -5089 172
rect -5181 132 -5089 138
rect -5023 172 -4931 178
rect -5023 138 -5011 172
rect -4943 138 -4931 172
rect -5023 132 -4931 138
rect -4865 172 -4773 178
rect -4865 138 -4853 172
rect -4785 138 -4773 172
rect -4865 132 -4773 138
rect -4707 172 -4615 178
rect -4707 138 -4695 172
rect -4627 138 -4615 172
rect -4707 132 -4615 138
rect -4549 172 -4457 178
rect -4549 138 -4537 172
rect -4469 138 -4457 172
rect -4549 132 -4457 138
rect -4391 172 -4299 178
rect -4391 138 -4379 172
rect -4311 138 -4299 172
rect -4391 132 -4299 138
rect -4233 172 -4141 178
rect -4233 138 -4221 172
rect -4153 138 -4141 172
rect -4233 132 -4141 138
rect -4075 172 -3983 178
rect -4075 138 -4063 172
rect -3995 138 -3983 172
rect -4075 132 -3983 138
rect -3917 172 -3825 178
rect -3917 138 -3905 172
rect -3837 138 -3825 172
rect -3917 132 -3825 138
rect -3759 172 -3667 178
rect -3759 138 -3747 172
rect -3679 138 -3667 172
rect -3759 132 -3667 138
rect -3601 172 -3509 178
rect -3601 138 -3589 172
rect -3521 138 -3509 172
rect -3601 132 -3509 138
rect -3443 172 -3351 178
rect -3443 138 -3431 172
rect -3363 138 -3351 172
rect -3443 132 -3351 138
rect -3285 172 -3193 178
rect -3285 138 -3273 172
rect -3205 138 -3193 172
rect -3285 132 -3193 138
rect -3127 172 -3035 178
rect -3127 138 -3115 172
rect -3047 138 -3035 172
rect -3127 132 -3035 138
rect -2969 172 -2877 178
rect -2969 138 -2957 172
rect -2889 138 -2877 172
rect -2969 132 -2877 138
rect -2811 172 -2719 178
rect -2811 138 -2799 172
rect -2731 138 -2719 172
rect -2811 132 -2719 138
rect -2653 172 -2561 178
rect -2653 138 -2641 172
rect -2573 138 -2561 172
rect -2653 132 -2561 138
rect -2495 172 -2403 178
rect -2495 138 -2483 172
rect -2415 138 -2403 172
rect -2495 132 -2403 138
rect -2337 172 -2245 178
rect -2337 138 -2325 172
rect -2257 138 -2245 172
rect -2337 132 -2245 138
rect -2179 172 -2087 178
rect -2179 138 -2167 172
rect -2099 138 -2087 172
rect -2179 132 -2087 138
rect -2021 172 -1929 178
rect -2021 138 -2009 172
rect -1941 138 -1929 172
rect -2021 132 -1929 138
rect -1863 172 -1771 178
rect -1863 138 -1851 172
rect -1783 138 -1771 172
rect -1863 132 -1771 138
rect -1705 172 -1613 178
rect -1705 138 -1693 172
rect -1625 138 -1613 172
rect -1705 132 -1613 138
rect -1547 172 -1455 178
rect -1547 138 -1535 172
rect -1467 138 -1455 172
rect -1547 132 -1455 138
rect -1389 172 -1297 178
rect -1389 138 -1377 172
rect -1309 138 -1297 172
rect -1389 132 -1297 138
rect -1231 172 -1139 178
rect -1231 138 -1219 172
rect -1151 138 -1139 172
rect -1231 132 -1139 138
rect -1073 172 -981 178
rect -1073 138 -1061 172
rect -993 138 -981 172
rect -1073 132 -981 138
rect -915 172 -823 178
rect -915 138 -903 172
rect -835 138 -823 172
rect -915 132 -823 138
rect -757 172 -665 178
rect -757 138 -745 172
rect -677 138 -665 172
rect -757 132 -665 138
rect -599 172 -507 178
rect -599 138 -587 172
rect -519 138 -507 172
rect -599 132 -507 138
rect -441 172 -349 178
rect -441 138 -429 172
rect -361 138 -349 172
rect -441 132 -349 138
rect -283 172 -191 178
rect -283 138 -271 172
rect -203 138 -191 172
rect -283 132 -191 138
rect -125 172 -33 178
rect -125 138 -113 172
rect -45 138 -33 172
rect -125 132 -33 138
rect 33 172 125 178
rect 33 138 45 172
rect 113 138 125 172
rect 33 132 125 138
rect 191 172 283 178
rect 191 138 203 172
rect 271 138 283 172
rect 191 132 283 138
rect 349 172 441 178
rect 349 138 361 172
rect 429 138 441 172
rect 349 132 441 138
rect 507 172 599 178
rect 507 138 519 172
rect 587 138 599 172
rect 507 132 599 138
rect 665 172 757 178
rect 665 138 677 172
rect 745 138 757 172
rect 665 132 757 138
rect 823 172 915 178
rect 823 138 835 172
rect 903 138 915 172
rect 823 132 915 138
rect 981 172 1073 178
rect 981 138 993 172
rect 1061 138 1073 172
rect 981 132 1073 138
rect 1139 172 1231 178
rect 1139 138 1151 172
rect 1219 138 1231 172
rect 1139 132 1231 138
rect 1297 172 1389 178
rect 1297 138 1309 172
rect 1377 138 1389 172
rect 1297 132 1389 138
rect 1455 172 1547 178
rect 1455 138 1467 172
rect 1535 138 1547 172
rect 1455 132 1547 138
rect 1613 172 1705 178
rect 1613 138 1625 172
rect 1693 138 1705 172
rect 1613 132 1705 138
rect 1771 172 1863 178
rect 1771 138 1783 172
rect 1851 138 1863 172
rect 1771 132 1863 138
rect 1929 172 2021 178
rect 1929 138 1941 172
rect 2009 138 2021 172
rect 1929 132 2021 138
rect 2087 172 2179 178
rect 2087 138 2099 172
rect 2167 138 2179 172
rect 2087 132 2179 138
rect 2245 172 2337 178
rect 2245 138 2257 172
rect 2325 138 2337 172
rect 2245 132 2337 138
rect 2403 172 2495 178
rect 2403 138 2415 172
rect 2483 138 2495 172
rect 2403 132 2495 138
rect 2561 172 2653 178
rect 2561 138 2573 172
rect 2641 138 2653 172
rect 2561 132 2653 138
rect 2719 172 2811 178
rect 2719 138 2731 172
rect 2799 138 2811 172
rect 2719 132 2811 138
rect 2877 172 2969 178
rect 2877 138 2889 172
rect 2957 138 2969 172
rect 2877 132 2969 138
rect 3035 172 3127 178
rect 3035 138 3047 172
rect 3115 138 3127 172
rect 3035 132 3127 138
rect 3193 172 3285 178
rect 3193 138 3205 172
rect 3273 138 3285 172
rect 3193 132 3285 138
rect 3351 172 3443 178
rect 3351 138 3363 172
rect 3431 138 3443 172
rect 3351 132 3443 138
rect 3509 172 3601 178
rect 3509 138 3521 172
rect 3589 138 3601 172
rect 3509 132 3601 138
rect 3667 172 3759 178
rect 3667 138 3679 172
rect 3747 138 3759 172
rect 3667 132 3759 138
rect 3825 172 3917 178
rect 3825 138 3837 172
rect 3905 138 3917 172
rect 3825 132 3917 138
rect 3983 172 4075 178
rect 3983 138 3995 172
rect 4063 138 4075 172
rect 3983 132 4075 138
rect 4141 172 4233 178
rect 4141 138 4153 172
rect 4221 138 4233 172
rect 4141 132 4233 138
rect 4299 172 4391 178
rect 4299 138 4311 172
rect 4379 138 4391 172
rect 4299 132 4391 138
rect 4457 172 4549 178
rect 4457 138 4469 172
rect 4537 138 4549 172
rect 4457 132 4549 138
rect 4615 172 4707 178
rect 4615 138 4627 172
rect 4695 138 4707 172
rect 4615 132 4707 138
rect 4773 172 4865 178
rect 4773 138 4785 172
rect 4853 138 4865 172
rect 4773 132 4865 138
rect 4931 172 5023 178
rect 4931 138 4943 172
rect 5011 138 5023 172
rect 4931 132 5023 138
rect 5089 172 5181 178
rect 5089 138 5101 172
rect 5169 138 5181 172
rect 5089 132 5181 138
rect 5247 172 5339 178
rect 5247 138 5259 172
rect 5327 138 5339 172
rect 5247 132 5339 138
rect 5405 172 5497 178
rect 5405 138 5417 172
rect 5485 138 5497 172
rect 5405 132 5497 138
rect 5563 172 5655 178
rect 5563 138 5575 172
rect 5643 138 5655 172
rect 5563 132 5655 138
rect 5721 172 5813 178
rect 5721 138 5733 172
rect 5801 138 5813 172
rect 5721 132 5813 138
rect 5879 172 5971 178
rect 5879 138 5891 172
rect 5959 138 5971 172
rect 5879 132 5971 138
rect 6037 172 6129 178
rect 6037 138 6049 172
rect 6117 138 6129 172
rect 6037 132 6129 138
rect 6195 172 6287 178
rect 6195 138 6207 172
rect 6275 138 6287 172
rect 6195 132 6287 138
rect 6353 172 6445 178
rect 6353 138 6365 172
rect 6433 138 6445 172
rect 6353 132 6445 138
rect 6511 172 6603 178
rect 6511 138 6523 172
rect 6591 138 6603 172
rect 6511 132 6603 138
rect 6669 172 6761 178
rect 6669 138 6681 172
rect 6749 138 6761 172
rect 6669 132 6761 138
rect 6827 172 6919 178
rect 6827 138 6839 172
rect 6907 138 6919 172
rect 6827 132 6919 138
rect 6985 172 7077 178
rect 6985 138 6997 172
rect 7065 138 7077 172
rect 6985 132 7077 138
rect 7143 172 7235 178
rect 7143 138 7155 172
rect 7223 138 7235 172
rect 7143 132 7235 138
rect 7301 172 7393 178
rect 7301 138 7313 172
rect 7381 138 7393 172
rect 7301 132 7393 138
rect 7459 172 7551 178
rect 7459 138 7471 172
rect 7539 138 7551 172
rect 7459 132 7551 138
rect 7617 172 7709 178
rect 7617 138 7629 172
rect 7697 138 7709 172
rect 7617 132 7709 138
rect 7775 172 7867 178
rect 7775 138 7787 172
rect 7855 138 7867 172
rect 7775 132 7867 138
rect 7933 172 8025 178
rect 7933 138 7945 172
rect 8013 138 8025 172
rect 7933 132 8025 138
rect 8091 172 8183 178
rect 8091 138 8103 172
rect 8171 138 8183 172
rect 8091 132 8183 138
rect 8249 172 8341 178
rect 8249 138 8261 172
rect 8329 138 8341 172
rect 8249 132 8341 138
rect 8407 172 8499 178
rect 8407 138 8419 172
rect 8487 138 8499 172
rect 8407 132 8499 138
rect 8565 172 8657 178
rect 8565 138 8577 172
rect 8645 138 8657 172
rect 8565 132 8657 138
rect 8723 172 8815 178
rect 8723 138 8735 172
rect 8803 138 8815 172
rect 8723 132 8815 138
rect 8881 172 8973 178
rect 8881 138 8893 172
rect 8961 138 8973 172
rect 8881 132 8973 138
rect 9039 172 9131 178
rect 9039 138 9051 172
rect 9119 138 9131 172
rect 9039 132 9131 138
rect 9197 172 9289 178
rect 9197 138 9209 172
rect 9277 138 9289 172
rect 9197 132 9289 138
rect 9355 172 9447 178
rect 9355 138 9367 172
rect 9435 138 9447 172
rect 9355 132 9447 138
rect -9503 88 -9457 100
rect -9503 -88 -9497 88
rect -9463 -88 -9457 88
rect -9503 -100 -9457 -88
rect -9345 88 -9299 100
rect -9345 -88 -9339 88
rect -9305 -88 -9299 88
rect -9345 -100 -9299 -88
rect -9187 88 -9141 100
rect -9187 -88 -9181 88
rect -9147 -88 -9141 88
rect -9187 -100 -9141 -88
rect -9029 88 -8983 100
rect -9029 -88 -9023 88
rect -8989 -88 -8983 88
rect -9029 -100 -8983 -88
rect -8871 88 -8825 100
rect -8871 -88 -8865 88
rect -8831 -88 -8825 88
rect -8871 -100 -8825 -88
rect -8713 88 -8667 100
rect -8713 -88 -8707 88
rect -8673 -88 -8667 88
rect -8713 -100 -8667 -88
rect -8555 88 -8509 100
rect -8555 -88 -8549 88
rect -8515 -88 -8509 88
rect -8555 -100 -8509 -88
rect -8397 88 -8351 100
rect -8397 -88 -8391 88
rect -8357 -88 -8351 88
rect -8397 -100 -8351 -88
rect -8239 88 -8193 100
rect -8239 -88 -8233 88
rect -8199 -88 -8193 88
rect -8239 -100 -8193 -88
rect -8081 88 -8035 100
rect -8081 -88 -8075 88
rect -8041 -88 -8035 88
rect -8081 -100 -8035 -88
rect -7923 88 -7877 100
rect -7923 -88 -7917 88
rect -7883 -88 -7877 88
rect -7923 -100 -7877 -88
rect -7765 88 -7719 100
rect -7765 -88 -7759 88
rect -7725 -88 -7719 88
rect -7765 -100 -7719 -88
rect -7607 88 -7561 100
rect -7607 -88 -7601 88
rect -7567 -88 -7561 88
rect -7607 -100 -7561 -88
rect -7449 88 -7403 100
rect -7449 -88 -7443 88
rect -7409 -88 -7403 88
rect -7449 -100 -7403 -88
rect -7291 88 -7245 100
rect -7291 -88 -7285 88
rect -7251 -88 -7245 88
rect -7291 -100 -7245 -88
rect -7133 88 -7087 100
rect -7133 -88 -7127 88
rect -7093 -88 -7087 88
rect -7133 -100 -7087 -88
rect -6975 88 -6929 100
rect -6975 -88 -6969 88
rect -6935 -88 -6929 88
rect -6975 -100 -6929 -88
rect -6817 88 -6771 100
rect -6817 -88 -6811 88
rect -6777 -88 -6771 88
rect -6817 -100 -6771 -88
rect -6659 88 -6613 100
rect -6659 -88 -6653 88
rect -6619 -88 -6613 88
rect -6659 -100 -6613 -88
rect -6501 88 -6455 100
rect -6501 -88 -6495 88
rect -6461 -88 -6455 88
rect -6501 -100 -6455 -88
rect -6343 88 -6297 100
rect -6343 -88 -6337 88
rect -6303 -88 -6297 88
rect -6343 -100 -6297 -88
rect -6185 88 -6139 100
rect -6185 -88 -6179 88
rect -6145 -88 -6139 88
rect -6185 -100 -6139 -88
rect -6027 88 -5981 100
rect -6027 -88 -6021 88
rect -5987 -88 -5981 88
rect -6027 -100 -5981 -88
rect -5869 88 -5823 100
rect -5869 -88 -5863 88
rect -5829 -88 -5823 88
rect -5869 -100 -5823 -88
rect -5711 88 -5665 100
rect -5711 -88 -5705 88
rect -5671 -88 -5665 88
rect -5711 -100 -5665 -88
rect -5553 88 -5507 100
rect -5553 -88 -5547 88
rect -5513 -88 -5507 88
rect -5553 -100 -5507 -88
rect -5395 88 -5349 100
rect -5395 -88 -5389 88
rect -5355 -88 -5349 88
rect -5395 -100 -5349 -88
rect -5237 88 -5191 100
rect -5237 -88 -5231 88
rect -5197 -88 -5191 88
rect -5237 -100 -5191 -88
rect -5079 88 -5033 100
rect -5079 -88 -5073 88
rect -5039 -88 -5033 88
rect -5079 -100 -5033 -88
rect -4921 88 -4875 100
rect -4921 -88 -4915 88
rect -4881 -88 -4875 88
rect -4921 -100 -4875 -88
rect -4763 88 -4717 100
rect -4763 -88 -4757 88
rect -4723 -88 -4717 88
rect -4763 -100 -4717 -88
rect -4605 88 -4559 100
rect -4605 -88 -4599 88
rect -4565 -88 -4559 88
rect -4605 -100 -4559 -88
rect -4447 88 -4401 100
rect -4447 -88 -4441 88
rect -4407 -88 -4401 88
rect -4447 -100 -4401 -88
rect -4289 88 -4243 100
rect -4289 -88 -4283 88
rect -4249 -88 -4243 88
rect -4289 -100 -4243 -88
rect -4131 88 -4085 100
rect -4131 -88 -4125 88
rect -4091 -88 -4085 88
rect -4131 -100 -4085 -88
rect -3973 88 -3927 100
rect -3973 -88 -3967 88
rect -3933 -88 -3927 88
rect -3973 -100 -3927 -88
rect -3815 88 -3769 100
rect -3815 -88 -3809 88
rect -3775 -88 -3769 88
rect -3815 -100 -3769 -88
rect -3657 88 -3611 100
rect -3657 -88 -3651 88
rect -3617 -88 -3611 88
rect -3657 -100 -3611 -88
rect -3499 88 -3453 100
rect -3499 -88 -3493 88
rect -3459 -88 -3453 88
rect -3499 -100 -3453 -88
rect -3341 88 -3295 100
rect -3341 -88 -3335 88
rect -3301 -88 -3295 88
rect -3341 -100 -3295 -88
rect -3183 88 -3137 100
rect -3183 -88 -3177 88
rect -3143 -88 -3137 88
rect -3183 -100 -3137 -88
rect -3025 88 -2979 100
rect -3025 -88 -3019 88
rect -2985 -88 -2979 88
rect -3025 -100 -2979 -88
rect -2867 88 -2821 100
rect -2867 -88 -2861 88
rect -2827 -88 -2821 88
rect -2867 -100 -2821 -88
rect -2709 88 -2663 100
rect -2709 -88 -2703 88
rect -2669 -88 -2663 88
rect -2709 -100 -2663 -88
rect -2551 88 -2505 100
rect -2551 -88 -2545 88
rect -2511 -88 -2505 88
rect -2551 -100 -2505 -88
rect -2393 88 -2347 100
rect -2393 -88 -2387 88
rect -2353 -88 -2347 88
rect -2393 -100 -2347 -88
rect -2235 88 -2189 100
rect -2235 -88 -2229 88
rect -2195 -88 -2189 88
rect -2235 -100 -2189 -88
rect -2077 88 -2031 100
rect -2077 -88 -2071 88
rect -2037 -88 -2031 88
rect -2077 -100 -2031 -88
rect -1919 88 -1873 100
rect -1919 -88 -1913 88
rect -1879 -88 -1873 88
rect -1919 -100 -1873 -88
rect -1761 88 -1715 100
rect -1761 -88 -1755 88
rect -1721 -88 -1715 88
rect -1761 -100 -1715 -88
rect -1603 88 -1557 100
rect -1603 -88 -1597 88
rect -1563 -88 -1557 88
rect -1603 -100 -1557 -88
rect -1445 88 -1399 100
rect -1445 -88 -1439 88
rect -1405 -88 -1399 88
rect -1445 -100 -1399 -88
rect -1287 88 -1241 100
rect -1287 -88 -1281 88
rect -1247 -88 -1241 88
rect -1287 -100 -1241 -88
rect -1129 88 -1083 100
rect -1129 -88 -1123 88
rect -1089 -88 -1083 88
rect -1129 -100 -1083 -88
rect -971 88 -925 100
rect -971 -88 -965 88
rect -931 -88 -925 88
rect -971 -100 -925 -88
rect -813 88 -767 100
rect -813 -88 -807 88
rect -773 -88 -767 88
rect -813 -100 -767 -88
rect -655 88 -609 100
rect -655 -88 -649 88
rect -615 -88 -609 88
rect -655 -100 -609 -88
rect -497 88 -451 100
rect -497 -88 -491 88
rect -457 -88 -451 88
rect -497 -100 -451 -88
rect -339 88 -293 100
rect -339 -88 -333 88
rect -299 -88 -293 88
rect -339 -100 -293 -88
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect 293 88 339 100
rect 293 -88 299 88
rect 333 -88 339 88
rect 293 -100 339 -88
rect 451 88 497 100
rect 451 -88 457 88
rect 491 -88 497 88
rect 451 -100 497 -88
rect 609 88 655 100
rect 609 -88 615 88
rect 649 -88 655 88
rect 609 -100 655 -88
rect 767 88 813 100
rect 767 -88 773 88
rect 807 -88 813 88
rect 767 -100 813 -88
rect 925 88 971 100
rect 925 -88 931 88
rect 965 -88 971 88
rect 925 -100 971 -88
rect 1083 88 1129 100
rect 1083 -88 1089 88
rect 1123 -88 1129 88
rect 1083 -100 1129 -88
rect 1241 88 1287 100
rect 1241 -88 1247 88
rect 1281 -88 1287 88
rect 1241 -100 1287 -88
rect 1399 88 1445 100
rect 1399 -88 1405 88
rect 1439 -88 1445 88
rect 1399 -100 1445 -88
rect 1557 88 1603 100
rect 1557 -88 1563 88
rect 1597 -88 1603 88
rect 1557 -100 1603 -88
rect 1715 88 1761 100
rect 1715 -88 1721 88
rect 1755 -88 1761 88
rect 1715 -100 1761 -88
rect 1873 88 1919 100
rect 1873 -88 1879 88
rect 1913 -88 1919 88
rect 1873 -100 1919 -88
rect 2031 88 2077 100
rect 2031 -88 2037 88
rect 2071 -88 2077 88
rect 2031 -100 2077 -88
rect 2189 88 2235 100
rect 2189 -88 2195 88
rect 2229 -88 2235 88
rect 2189 -100 2235 -88
rect 2347 88 2393 100
rect 2347 -88 2353 88
rect 2387 -88 2393 88
rect 2347 -100 2393 -88
rect 2505 88 2551 100
rect 2505 -88 2511 88
rect 2545 -88 2551 88
rect 2505 -100 2551 -88
rect 2663 88 2709 100
rect 2663 -88 2669 88
rect 2703 -88 2709 88
rect 2663 -100 2709 -88
rect 2821 88 2867 100
rect 2821 -88 2827 88
rect 2861 -88 2867 88
rect 2821 -100 2867 -88
rect 2979 88 3025 100
rect 2979 -88 2985 88
rect 3019 -88 3025 88
rect 2979 -100 3025 -88
rect 3137 88 3183 100
rect 3137 -88 3143 88
rect 3177 -88 3183 88
rect 3137 -100 3183 -88
rect 3295 88 3341 100
rect 3295 -88 3301 88
rect 3335 -88 3341 88
rect 3295 -100 3341 -88
rect 3453 88 3499 100
rect 3453 -88 3459 88
rect 3493 -88 3499 88
rect 3453 -100 3499 -88
rect 3611 88 3657 100
rect 3611 -88 3617 88
rect 3651 -88 3657 88
rect 3611 -100 3657 -88
rect 3769 88 3815 100
rect 3769 -88 3775 88
rect 3809 -88 3815 88
rect 3769 -100 3815 -88
rect 3927 88 3973 100
rect 3927 -88 3933 88
rect 3967 -88 3973 88
rect 3927 -100 3973 -88
rect 4085 88 4131 100
rect 4085 -88 4091 88
rect 4125 -88 4131 88
rect 4085 -100 4131 -88
rect 4243 88 4289 100
rect 4243 -88 4249 88
rect 4283 -88 4289 88
rect 4243 -100 4289 -88
rect 4401 88 4447 100
rect 4401 -88 4407 88
rect 4441 -88 4447 88
rect 4401 -100 4447 -88
rect 4559 88 4605 100
rect 4559 -88 4565 88
rect 4599 -88 4605 88
rect 4559 -100 4605 -88
rect 4717 88 4763 100
rect 4717 -88 4723 88
rect 4757 -88 4763 88
rect 4717 -100 4763 -88
rect 4875 88 4921 100
rect 4875 -88 4881 88
rect 4915 -88 4921 88
rect 4875 -100 4921 -88
rect 5033 88 5079 100
rect 5033 -88 5039 88
rect 5073 -88 5079 88
rect 5033 -100 5079 -88
rect 5191 88 5237 100
rect 5191 -88 5197 88
rect 5231 -88 5237 88
rect 5191 -100 5237 -88
rect 5349 88 5395 100
rect 5349 -88 5355 88
rect 5389 -88 5395 88
rect 5349 -100 5395 -88
rect 5507 88 5553 100
rect 5507 -88 5513 88
rect 5547 -88 5553 88
rect 5507 -100 5553 -88
rect 5665 88 5711 100
rect 5665 -88 5671 88
rect 5705 -88 5711 88
rect 5665 -100 5711 -88
rect 5823 88 5869 100
rect 5823 -88 5829 88
rect 5863 -88 5869 88
rect 5823 -100 5869 -88
rect 5981 88 6027 100
rect 5981 -88 5987 88
rect 6021 -88 6027 88
rect 5981 -100 6027 -88
rect 6139 88 6185 100
rect 6139 -88 6145 88
rect 6179 -88 6185 88
rect 6139 -100 6185 -88
rect 6297 88 6343 100
rect 6297 -88 6303 88
rect 6337 -88 6343 88
rect 6297 -100 6343 -88
rect 6455 88 6501 100
rect 6455 -88 6461 88
rect 6495 -88 6501 88
rect 6455 -100 6501 -88
rect 6613 88 6659 100
rect 6613 -88 6619 88
rect 6653 -88 6659 88
rect 6613 -100 6659 -88
rect 6771 88 6817 100
rect 6771 -88 6777 88
rect 6811 -88 6817 88
rect 6771 -100 6817 -88
rect 6929 88 6975 100
rect 6929 -88 6935 88
rect 6969 -88 6975 88
rect 6929 -100 6975 -88
rect 7087 88 7133 100
rect 7087 -88 7093 88
rect 7127 -88 7133 88
rect 7087 -100 7133 -88
rect 7245 88 7291 100
rect 7245 -88 7251 88
rect 7285 -88 7291 88
rect 7245 -100 7291 -88
rect 7403 88 7449 100
rect 7403 -88 7409 88
rect 7443 -88 7449 88
rect 7403 -100 7449 -88
rect 7561 88 7607 100
rect 7561 -88 7567 88
rect 7601 -88 7607 88
rect 7561 -100 7607 -88
rect 7719 88 7765 100
rect 7719 -88 7725 88
rect 7759 -88 7765 88
rect 7719 -100 7765 -88
rect 7877 88 7923 100
rect 7877 -88 7883 88
rect 7917 -88 7923 88
rect 7877 -100 7923 -88
rect 8035 88 8081 100
rect 8035 -88 8041 88
rect 8075 -88 8081 88
rect 8035 -100 8081 -88
rect 8193 88 8239 100
rect 8193 -88 8199 88
rect 8233 -88 8239 88
rect 8193 -100 8239 -88
rect 8351 88 8397 100
rect 8351 -88 8357 88
rect 8391 -88 8397 88
rect 8351 -100 8397 -88
rect 8509 88 8555 100
rect 8509 -88 8515 88
rect 8549 -88 8555 88
rect 8509 -100 8555 -88
rect 8667 88 8713 100
rect 8667 -88 8673 88
rect 8707 -88 8713 88
rect 8667 -100 8713 -88
rect 8825 88 8871 100
rect 8825 -88 8831 88
rect 8865 -88 8871 88
rect 8825 -100 8871 -88
rect 8983 88 9029 100
rect 8983 -88 8989 88
rect 9023 -88 9029 88
rect 8983 -100 9029 -88
rect 9141 88 9187 100
rect 9141 -88 9147 88
rect 9181 -88 9187 88
rect 9141 -100 9187 -88
rect 9299 88 9345 100
rect 9299 -88 9305 88
rect 9339 -88 9345 88
rect 9299 -100 9345 -88
rect 9457 88 9503 100
rect 9457 -88 9463 88
rect 9497 -88 9503 88
rect 9457 -100 9503 -88
rect -9447 -138 -9355 -132
rect -9447 -172 -9435 -138
rect -9367 -172 -9355 -138
rect -9447 -178 -9355 -172
rect -9289 -138 -9197 -132
rect -9289 -172 -9277 -138
rect -9209 -172 -9197 -138
rect -9289 -178 -9197 -172
rect -9131 -138 -9039 -132
rect -9131 -172 -9119 -138
rect -9051 -172 -9039 -138
rect -9131 -178 -9039 -172
rect -8973 -138 -8881 -132
rect -8973 -172 -8961 -138
rect -8893 -172 -8881 -138
rect -8973 -178 -8881 -172
rect -8815 -138 -8723 -132
rect -8815 -172 -8803 -138
rect -8735 -172 -8723 -138
rect -8815 -178 -8723 -172
rect -8657 -138 -8565 -132
rect -8657 -172 -8645 -138
rect -8577 -172 -8565 -138
rect -8657 -178 -8565 -172
rect -8499 -138 -8407 -132
rect -8499 -172 -8487 -138
rect -8419 -172 -8407 -138
rect -8499 -178 -8407 -172
rect -8341 -138 -8249 -132
rect -8341 -172 -8329 -138
rect -8261 -172 -8249 -138
rect -8341 -178 -8249 -172
rect -8183 -138 -8091 -132
rect -8183 -172 -8171 -138
rect -8103 -172 -8091 -138
rect -8183 -178 -8091 -172
rect -8025 -138 -7933 -132
rect -8025 -172 -8013 -138
rect -7945 -172 -7933 -138
rect -8025 -178 -7933 -172
rect -7867 -138 -7775 -132
rect -7867 -172 -7855 -138
rect -7787 -172 -7775 -138
rect -7867 -178 -7775 -172
rect -7709 -138 -7617 -132
rect -7709 -172 -7697 -138
rect -7629 -172 -7617 -138
rect -7709 -178 -7617 -172
rect -7551 -138 -7459 -132
rect -7551 -172 -7539 -138
rect -7471 -172 -7459 -138
rect -7551 -178 -7459 -172
rect -7393 -138 -7301 -132
rect -7393 -172 -7381 -138
rect -7313 -172 -7301 -138
rect -7393 -178 -7301 -172
rect -7235 -138 -7143 -132
rect -7235 -172 -7223 -138
rect -7155 -172 -7143 -138
rect -7235 -178 -7143 -172
rect -7077 -138 -6985 -132
rect -7077 -172 -7065 -138
rect -6997 -172 -6985 -138
rect -7077 -178 -6985 -172
rect -6919 -138 -6827 -132
rect -6919 -172 -6907 -138
rect -6839 -172 -6827 -138
rect -6919 -178 -6827 -172
rect -6761 -138 -6669 -132
rect -6761 -172 -6749 -138
rect -6681 -172 -6669 -138
rect -6761 -178 -6669 -172
rect -6603 -138 -6511 -132
rect -6603 -172 -6591 -138
rect -6523 -172 -6511 -138
rect -6603 -178 -6511 -172
rect -6445 -138 -6353 -132
rect -6445 -172 -6433 -138
rect -6365 -172 -6353 -138
rect -6445 -178 -6353 -172
rect -6287 -138 -6195 -132
rect -6287 -172 -6275 -138
rect -6207 -172 -6195 -138
rect -6287 -178 -6195 -172
rect -6129 -138 -6037 -132
rect -6129 -172 -6117 -138
rect -6049 -172 -6037 -138
rect -6129 -178 -6037 -172
rect -5971 -138 -5879 -132
rect -5971 -172 -5959 -138
rect -5891 -172 -5879 -138
rect -5971 -178 -5879 -172
rect -5813 -138 -5721 -132
rect -5813 -172 -5801 -138
rect -5733 -172 -5721 -138
rect -5813 -178 -5721 -172
rect -5655 -138 -5563 -132
rect -5655 -172 -5643 -138
rect -5575 -172 -5563 -138
rect -5655 -178 -5563 -172
rect -5497 -138 -5405 -132
rect -5497 -172 -5485 -138
rect -5417 -172 -5405 -138
rect -5497 -178 -5405 -172
rect -5339 -138 -5247 -132
rect -5339 -172 -5327 -138
rect -5259 -172 -5247 -138
rect -5339 -178 -5247 -172
rect -5181 -138 -5089 -132
rect -5181 -172 -5169 -138
rect -5101 -172 -5089 -138
rect -5181 -178 -5089 -172
rect -5023 -138 -4931 -132
rect -5023 -172 -5011 -138
rect -4943 -172 -4931 -138
rect -5023 -178 -4931 -172
rect -4865 -138 -4773 -132
rect -4865 -172 -4853 -138
rect -4785 -172 -4773 -138
rect -4865 -178 -4773 -172
rect -4707 -138 -4615 -132
rect -4707 -172 -4695 -138
rect -4627 -172 -4615 -138
rect -4707 -178 -4615 -172
rect -4549 -138 -4457 -132
rect -4549 -172 -4537 -138
rect -4469 -172 -4457 -138
rect -4549 -178 -4457 -172
rect -4391 -138 -4299 -132
rect -4391 -172 -4379 -138
rect -4311 -172 -4299 -138
rect -4391 -178 -4299 -172
rect -4233 -138 -4141 -132
rect -4233 -172 -4221 -138
rect -4153 -172 -4141 -138
rect -4233 -178 -4141 -172
rect -4075 -138 -3983 -132
rect -4075 -172 -4063 -138
rect -3995 -172 -3983 -138
rect -4075 -178 -3983 -172
rect -3917 -138 -3825 -132
rect -3917 -172 -3905 -138
rect -3837 -172 -3825 -138
rect -3917 -178 -3825 -172
rect -3759 -138 -3667 -132
rect -3759 -172 -3747 -138
rect -3679 -172 -3667 -138
rect -3759 -178 -3667 -172
rect -3601 -138 -3509 -132
rect -3601 -172 -3589 -138
rect -3521 -172 -3509 -138
rect -3601 -178 -3509 -172
rect -3443 -138 -3351 -132
rect -3443 -172 -3431 -138
rect -3363 -172 -3351 -138
rect -3443 -178 -3351 -172
rect -3285 -138 -3193 -132
rect -3285 -172 -3273 -138
rect -3205 -172 -3193 -138
rect -3285 -178 -3193 -172
rect -3127 -138 -3035 -132
rect -3127 -172 -3115 -138
rect -3047 -172 -3035 -138
rect -3127 -178 -3035 -172
rect -2969 -138 -2877 -132
rect -2969 -172 -2957 -138
rect -2889 -172 -2877 -138
rect -2969 -178 -2877 -172
rect -2811 -138 -2719 -132
rect -2811 -172 -2799 -138
rect -2731 -172 -2719 -138
rect -2811 -178 -2719 -172
rect -2653 -138 -2561 -132
rect -2653 -172 -2641 -138
rect -2573 -172 -2561 -138
rect -2653 -178 -2561 -172
rect -2495 -138 -2403 -132
rect -2495 -172 -2483 -138
rect -2415 -172 -2403 -138
rect -2495 -178 -2403 -172
rect -2337 -138 -2245 -132
rect -2337 -172 -2325 -138
rect -2257 -172 -2245 -138
rect -2337 -178 -2245 -172
rect -2179 -138 -2087 -132
rect -2179 -172 -2167 -138
rect -2099 -172 -2087 -138
rect -2179 -178 -2087 -172
rect -2021 -138 -1929 -132
rect -2021 -172 -2009 -138
rect -1941 -172 -1929 -138
rect -2021 -178 -1929 -172
rect -1863 -138 -1771 -132
rect -1863 -172 -1851 -138
rect -1783 -172 -1771 -138
rect -1863 -178 -1771 -172
rect -1705 -138 -1613 -132
rect -1705 -172 -1693 -138
rect -1625 -172 -1613 -138
rect -1705 -178 -1613 -172
rect -1547 -138 -1455 -132
rect -1547 -172 -1535 -138
rect -1467 -172 -1455 -138
rect -1547 -178 -1455 -172
rect -1389 -138 -1297 -132
rect -1389 -172 -1377 -138
rect -1309 -172 -1297 -138
rect -1389 -178 -1297 -172
rect -1231 -138 -1139 -132
rect -1231 -172 -1219 -138
rect -1151 -172 -1139 -138
rect -1231 -178 -1139 -172
rect -1073 -138 -981 -132
rect -1073 -172 -1061 -138
rect -993 -172 -981 -138
rect -1073 -178 -981 -172
rect -915 -138 -823 -132
rect -915 -172 -903 -138
rect -835 -172 -823 -138
rect -915 -178 -823 -172
rect -757 -138 -665 -132
rect -757 -172 -745 -138
rect -677 -172 -665 -138
rect -757 -178 -665 -172
rect -599 -138 -507 -132
rect -599 -172 -587 -138
rect -519 -172 -507 -138
rect -599 -178 -507 -172
rect -441 -138 -349 -132
rect -441 -172 -429 -138
rect -361 -172 -349 -138
rect -441 -178 -349 -172
rect -283 -138 -191 -132
rect -283 -172 -271 -138
rect -203 -172 -191 -138
rect -283 -178 -191 -172
rect -125 -138 -33 -132
rect -125 -172 -113 -138
rect -45 -172 -33 -138
rect -125 -178 -33 -172
rect 33 -138 125 -132
rect 33 -172 45 -138
rect 113 -172 125 -138
rect 33 -178 125 -172
rect 191 -138 283 -132
rect 191 -172 203 -138
rect 271 -172 283 -138
rect 191 -178 283 -172
rect 349 -138 441 -132
rect 349 -172 361 -138
rect 429 -172 441 -138
rect 349 -178 441 -172
rect 507 -138 599 -132
rect 507 -172 519 -138
rect 587 -172 599 -138
rect 507 -178 599 -172
rect 665 -138 757 -132
rect 665 -172 677 -138
rect 745 -172 757 -138
rect 665 -178 757 -172
rect 823 -138 915 -132
rect 823 -172 835 -138
rect 903 -172 915 -138
rect 823 -178 915 -172
rect 981 -138 1073 -132
rect 981 -172 993 -138
rect 1061 -172 1073 -138
rect 981 -178 1073 -172
rect 1139 -138 1231 -132
rect 1139 -172 1151 -138
rect 1219 -172 1231 -138
rect 1139 -178 1231 -172
rect 1297 -138 1389 -132
rect 1297 -172 1309 -138
rect 1377 -172 1389 -138
rect 1297 -178 1389 -172
rect 1455 -138 1547 -132
rect 1455 -172 1467 -138
rect 1535 -172 1547 -138
rect 1455 -178 1547 -172
rect 1613 -138 1705 -132
rect 1613 -172 1625 -138
rect 1693 -172 1705 -138
rect 1613 -178 1705 -172
rect 1771 -138 1863 -132
rect 1771 -172 1783 -138
rect 1851 -172 1863 -138
rect 1771 -178 1863 -172
rect 1929 -138 2021 -132
rect 1929 -172 1941 -138
rect 2009 -172 2021 -138
rect 1929 -178 2021 -172
rect 2087 -138 2179 -132
rect 2087 -172 2099 -138
rect 2167 -172 2179 -138
rect 2087 -178 2179 -172
rect 2245 -138 2337 -132
rect 2245 -172 2257 -138
rect 2325 -172 2337 -138
rect 2245 -178 2337 -172
rect 2403 -138 2495 -132
rect 2403 -172 2415 -138
rect 2483 -172 2495 -138
rect 2403 -178 2495 -172
rect 2561 -138 2653 -132
rect 2561 -172 2573 -138
rect 2641 -172 2653 -138
rect 2561 -178 2653 -172
rect 2719 -138 2811 -132
rect 2719 -172 2731 -138
rect 2799 -172 2811 -138
rect 2719 -178 2811 -172
rect 2877 -138 2969 -132
rect 2877 -172 2889 -138
rect 2957 -172 2969 -138
rect 2877 -178 2969 -172
rect 3035 -138 3127 -132
rect 3035 -172 3047 -138
rect 3115 -172 3127 -138
rect 3035 -178 3127 -172
rect 3193 -138 3285 -132
rect 3193 -172 3205 -138
rect 3273 -172 3285 -138
rect 3193 -178 3285 -172
rect 3351 -138 3443 -132
rect 3351 -172 3363 -138
rect 3431 -172 3443 -138
rect 3351 -178 3443 -172
rect 3509 -138 3601 -132
rect 3509 -172 3521 -138
rect 3589 -172 3601 -138
rect 3509 -178 3601 -172
rect 3667 -138 3759 -132
rect 3667 -172 3679 -138
rect 3747 -172 3759 -138
rect 3667 -178 3759 -172
rect 3825 -138 3917 -132
rect 3825 -172 3837 -138
rect 3905 -172 3917 -138
rect 3825 -178 3917 -172
rect 3983 -138 4075 -132
rect 3983 -172 3995 -138
rect 4063 -172 4075 -138
rect 3983 -178 4075 -172
rect 4141 -138 4233 -132
rect 4141 -172 4153 -138
rect 4221 -172 4233 -138
rect 4141 -178 4233 -172
rect 4299 -138 4391 -132
rect 4299 -172 4311 -138
rect 4379 -172 4391 -138
rect 4299 -178 4391 -172
rect 4457 -138 4549 -132
rect 4457 -172 4469 -138
rect 4537 -172 4549 -138
rect 4457 -178 4549 -172
rect 4615 -138 4707 -132
rect 4615 -172 4627 -138
rect 4695 -172 4707 -138
rect 4615 -178 4707 -172
rect 4773 -138 4865 -132
rect 4773 -172 4785 -138
rect 4853 -172 4865 -138
rect 4773 -178 4865 -172
rect 4931 -138 5023 -132
rect 4931 -172 4943 -138
rect 5011 -172 5023 -138
rect 4931 -178 5023 -172
rect 5089 -138 5181 -132
rect 5089 -172 5101 -138
rect 5169 -172 5181 -138
rect 5089 -178 5181 -172
rect 5247 -138 5339 -132
rect 5247 -172 5259 -138
rect 5327 -172 5339 -138
rect 5247 -178 5339 -172
rect 5405 -138 5497 -132
rect 5405 -172 5417 -138
rect 5485 -172 5497 -138
rect 5405 -178 5497 -172
rect 5563 -138 5655 -132
rect 5563 -172 5575 -138
rect 5643 -172 5655 -138
rect 5563 -178 5655 -172
rect 5721 -138 5813 -132
rect 5721 -172 5733 -138
rect 5801 -172 5813 -138
rect 5721 -178 5813 -172
rect 5879 -138 5971 -132
rect 5879 -172 5891 -138
rect 5959 -172 5971 -138
rect 5879 -178 5971 -172
rect 6037 -138 6129 -132
rect 6037 -172 6049 -138
rect 6117 -172 6129 -138
rect 6037 -178 6129 -172
rect 6195 -138 6287 -132
rect 6195 -172 6207 -138
rect 6275 -172 6287 -138
rect 6195 -178 6287 -172
rect 6353 -138 6445 -132
rect 6353 -172 6365 -138
rect 6433 -172 6445 -138
rect 6353 -178 6445 -172
rect 6511 -138 6603 -132
rect 6511 -172 6523 -138
rect 6591 -172 6603 -138
rect 6511 -178 6603 -172
rect 6669 -138 6761 -132
rect 6669 -172 6681 -138
rect 6749 -172 6761 -138
rect 6669 -178 6761 -172
rect 6827 -138 6919 -132
rect 6827 -172 6839 -138
rect 6907 -172 6919 -138
rect 6827 -178 6919 -172
rect 6985 -138 7077 -132
rect 6985 -172 6997 -138
rect 7065 -172 7077 -138
rect 6985 -178 7077 -172
rect 7143 -138 7235 -132
rect 7143 -172 7155 -138
rect 7223 -172 7235 -138
rect 7143 -178 7235 -172
rect 7301 -138 7393 -132
rect 7301 -172 7313 -138
rect 7381 -172 7393 -138
rect 7301 -178 7393 -172
rect 7459 -138 7551 -132
rect 7459 -172 7471 -138
rect 7539 -172 7551 -138
rect 7459 -178 7551 -172
rect 7617 -138 7709 -132
rect 7617 -172 7629 -138
rect 7697 -172 7709 -138
rect 7617 -178 7709 -172
rect 7775 -138 7867 -132
rect 7775 -172 7787 -138
rect 7855 -172 7867 -138
rect 7775 -178 7867 -172
rect 7933 -138 8025 -132
rect 7933 -172 7945 -138
rect 8013 -172 8025 -138
rect 7933 -178 8025 -172
rect 8091 -138 8183 -132
rect 8091 -172 8103 -138
rect 8171 -172 8183 -138
rect 8091 -178 8183 -172
rect 8249 -138 8341 -132
rect 8249 -172 8261 -138
rect 8329 -172 8341 -138
rect 8249 -178 8341 -172
rect 8407 -138 8499 -132
rect 8407 -172 8419 -138
rect 8487 -172 8499 -138
rect 8407 -178 8499 -172
rect 8565 -138 8657 -132
rect 8565 -172 8577 -138
rect 8645 -172 8657 -138
rect 8565 -178 8657 -172
rect 8723 -138 8815 -132
rect 8723 -172 8735 -138
rect 8803 -172 8815 -138
rect 8723 -178 8815 -172
rect 8881 -138 8973 -132
rect 8881 -172 8893 -138
rect 8961 -172 8973 -138
rect 8881 -178 8973 -172
rect 9039 -138 9131 -132
rect 9039 -172 9051 -138
rect 9119 -172 9131 -138
rect 9039 -178 9131 -172
rect 9197 -138 9289 -132
rect 9197 -172 9209 -138
rect 9277 -172 9289 -138
rect 9197 -178 9289 -172
rect 9355 -138 9447 -132
rect 9355 -172 9367 -138
rect 9435 -172 9447 -138
rect 9355 -178 9447 -172
<< properties >>
string FIXED_BBOX -9614 -293 9614 293
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 120 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
