magic
tech sky130A
magscale 1 2
timestamp 1722642941
<< checkpaint >>
rect 73830 -17337 76752 -13553
<< error_s >>
rect -19917 -11529 -19900 -10913
rect -19863 -11583 -19846 -10962
rect -19336 -10974 -19221 -10962
rect -19329 -11008 -19221 -10974
rect -19336 -11020 -19221 -11008
rect -19279 -11075 -19221 -11020
rect -19238 -11212 -19221 -11075
rect -19845 -11690 -19289 -11328
rect -19279 -11566 -19221 -11212
rect -19238 -11624 -19221 -11566
rect -19220 -11075 -19155 -11039
rect -19220 -11133 -19069 -11075
rect -19220 -11624 -19126 -11133
rect -19220 -11690 -19155 -11624
rect -18747 -11677 -18700 -11375
rect -19141 -11699 -18700 -11677
rect -18693 -11699 -18646 -11429
rect -18559 -11677 -18534 -11674
rect -19141 -11707 -18712 -11699
rect -18681 -11711 -18678 -11699
rect -19107 -11741 -18678 -11711
rect -18559 -11745 -18525 -11677
rect -18559 -11767 -18527 -11749
rect -18559 -11783 -18511 -11767
rect -18501 -11771 -18499 -11685
rect -18401 -11767 -18369 -11749
rect -18563 -11799 -18511 -11783
rect -18693 -11867 -18646 -11802
rect -18642 -11849 -18635 -11802
rect -18577 -11813 -18511 -11799
rect -18501 -11813 -18469 -11791
rect -18401 -11813 -18353 -11767
rect -18343 -11813 -18311 -11791
rect -18577 -11819 -18311 -11813
rect -18589 -11833 -18311 -11819
rect -18611 -11851 -18311 -11833
rect -18273 -11826 -18243 -11797
rect -18231 -11826 -18197 -11817
rect -18273 -11827 -18197 -11826
rect -18185 -11827 -18147 -11791
rect -18273 -11851 -18147 -11827
rect -18693 -11921 -18635 -11867
rect -18595 -11883 -18588 -11851
rect -18585 -11855 -18453 -11851
rect -18451 -11855 -18295 -11851
rect -18585 -11875 -18295 -11855
rect -18585 -11877 -18249 -11875
rect -18559 -11917 -18249 -11877
rect -18559 -11921 -18407 -11917
rect -18401 -11921 -18249 -11917
rect -18219 -11889 -18173 -11851
rect -18769 -11933 -18635 -11921
rect -18611 -11933 -18575 -11921
rect -18501 -11923 -18379 -11921
rect -18343 -11923 -18243 -11921
rect -18219 -11923 -18212 -11889
rect -18501 -11933 -18407 -11923
rect -18353 -11933 -18243 -11923
rect -18185 -11928 -18173 -11889
rect -18161 -11923 -18114 -11892
rect -18693 -11955 -18575 -11933
rect -18511 -11939 -18439 -11933
rect -18353 -11939 -18223 -11933
rect -18185 -11939 -18150 -11928
rect -18511 -11940 -18452 -11939
rect -18511 -11955 -18453 -11940
rect -18353 -11955 -18281 -11939
rect -18693 -11959 -18281 -11955
rect -18693 -11965 -18511 -11959
rect -18693 -12015 -18635 -11965
rect -18623 -12013 -18511 -11965
rect -18501 -11961 -18465 -11959
rect -18501 -11993 -18485 -11961
rect -18501 -12005 -18465 -11993
rect -18499 -12013 -18465 -12005
rect -18453 -12013 -18353 -11959
rect -18343 -11961 -18307 -11959
rect -18343 -11993 -18327 -11961
rect -18343 -12005 -18307 -11993
rect -18341 -12013 -18307 -12005
rect -18623 -12015 -18295 -12013
rect -18693 -12019 -18623 -12015
rect -18611 -12019 -18586 -12015
rect -18536 -12019 -18511 -12015
rect -18499 -12019 -18465 -12015
rect -18453 -12019 -18428 -12015
rect -18378 -12019 -18353 -12015
rect -18341 -12019 -18307 -12015
rect -18693 -12039 -18299 -12019
rect -18295 -12039 -18270 -12015
rect -18693 -12040 -18270 -12039
rect -18693 -12048 -18273 -12040
rect -18693 -12061 -18270 -12048
rect -17750 -12061 -17747 -11441
rect -18693 -12063 -18299 -12061
rect -18295 -12063 -18270 -12061
rect -18693 -12073 -18270 -12063
rect -17716 -12073 -17682 -11375
rect -17420 -11733 -17386 -11647
rect -17445 -11799 -17350 -11733
rect -17445 -11857 -17234 -11799
rect 14432 -11811 14547 -11799
rect 14439 -11845 14547 -11811
rect 14432 -11857 14547 -11845
rect -18729 -12121 -18669 -12073
rect -18611 -12121 -18511 -12073
rect -18453 -12121 -18353 -12073
rect -17716 -12095 -17713 -12073
rect -18623 -12155 -18611 -12121
rect -18511 -12155 -18499 -12121
rect -18465 -12155 -18453 -12121
rect -18353 -12155 -18341 -12121
rect -18307 -12155 -18295 -12121
rect -17445 -12396 -17321 -11857
rect 14489 -11912 14547 -11857
rect -17245 -12230 -17234 -12030
rect -17445 -12432 -17350 -12396
rect 14530 -12461 14547 -11912
rect 14548 -11912 14613 -11876
rect 14548 -11970 14699 -11912
rect 14548 -12461 14642 -11970
rect 33230 -12338 33250 -12244
rect 33374 -12266 33408 -12244
rect 33532 -12266 33566 -12244
rect 33252 -12324 33736 -12266
rect 33252 -12340 33310 -12324
rect 33678 -12334 33736 -12324
rect 33678 -12338 33709 -12334
rect 33252 -12372 33332 -12340
rect 33678 -12372 33712 -12338
rect 33262 -12422 33310 -12372
rect 33436 -12382 33504 -12378
rect 33420 -12406 33520 -12382
rect 14548 -12527 14613 -12461
rect 33264 -12510 33298 -12422
rect 33444 -12440 33544 -12416
rect 33578 -12422 33586 -12372
rect 33656 -12374 33712 -12372
rect 33656 -12406 33724 -12374
rect 33678 -12422 33689 -12406
rect 33460 -12444 33528 -12440
rect 33398 -12498 33432 -12484
rect 33556 -12498 33590 -12484
rect 33386 -12510 33602 -12498
rect 33690 -12510 33724 -12406
rect 31956 -12544 33762 -12510
rect 33264 -12802 33298 -12544
rect 33386 -12556 33602 -12544
rect 33690 -12802 33724 -12544
rect 33823 -12556 33870 -11923
rect 33877 -12610 33924 -11977
rect 34303 -12247 34361 -12161
rect 34302 -12313 34397 -12247
rect 34302 -12371 34513 -12313
rect 34302 -12621 34426 -12371
rect 34502 -12621 34513 -12544
rect 34302 -12657 34415 -12621
rect 34368 -12675 34415 -12657
rect 34835 -12975 34852 -12359
rect 34889 -13024 34906 -12408
rect 35514 -13070 35531 -12454
rect 35568 -13119 35585 -12503
rect 36193 -13165 36210 -12549
rect 36247 -13219 36264 -12598
rect 36774 -12610 36889 -12598
rect 36781 -12644 36889 -12610
rect 36774 -12656 36889 -12644
rect 36831 -12711 36889 -12656
rect 36872 -12848 36889 -12711
rect 36265 -13202 36821 -12964
rect 36831 -13202 36889 -12848
rect 36265 -13260 36889 -13202
rect 36890 -12711 36955 -12675
rect 36890 -12769 37041 -12711
rect 36890 -13260 36984 -12769
rect 36265 -13318 36821 -13260
rect 36890 -13318 36955 -13260
rect 36265 -13326 36955 -13318
rect 36738 -13644 36785 -13326
rect 36938 -13343 37298 -13332
rect 36792 -13698 36839 -13354
rect 37363 -13355 37410 -13011
rect 36904 -13377 37264 -13366
rect 37417 -13409 37464 -13065
rect 37229 -13998 37276 -13654
rect 37429 -13697 37789 -13686
rect 37283 -14052 37330 -13708
rect 37854 -13709 37901 -13365
rect 37395 -13731 37755 -13720
rect 37908 -13763 37955 -13419
rect 37720 -14352 37767 -14008
rect 37920 -14051 38280 -14040
rect 37774 -14406 37821 -14062
rect 38345 -14063 38392 -13719
rect 37886 -14085 38246 -14074
rect 38399 -14117 38446 -13773
rect 38825 -14043 38883 -13957
rect 38824 -14109 38919 -14043
rect 38824 -14167 39035 -14109
rect 38824 -14417 38948 -14167
rect 39024 -14417 39035 -14340
rect 38824 -14453 38937 -14417
rect 38890 -14471 38937 -14453
rect 39515 -14771 39532 -14155
rect 39569 -14825 39586 -14204
rect 40096 -14216 40211 -14204
rect 40103 -14250 40211 -14216
rect 40096 -14262 40211 -14250
rect 40153 -14317 40211 -14262
rect 40194 -14454 40211 -14317
rect 39587 -14932 40143 -14570
rect 40153 -14808 40211 -14454
rect 40194 -14866 40211 -14808
rect 40212 -14317 40277 -14281
rect 40212 -14375 40363 -14317
rect 40212 -14866 40306 -14375
rect 40212 -14932 40277 -14866
rect 40685 -14961 40732 -14617
rect 40739 -15015 40786 -14671
rect 41176 -15315 41223 -14682
rect 41655 -14736 41750 -14717
rect 41230 -15369 41277 -14736
rect 41569 -14783 41750 -14736
rect 41655 -14841 41866 -14783
rect 41655 -15380 41779 -14841
rect 41855 -15214 41866 -15014
rect 73455 -15202 73513 -15086
rect 73589 -15202 73647 -15082
rect 73660 -15202 73713 -15198
rect 73336 -15234 73713 -15202
rect 73336 -15238 73799 -15234
rect 73336 -15268 73856 -15238
rect 73336 -15372 73730 -15268
rect 73798 -15336 73799 -15296
rect 73810 -15336 73844 -15314
rect 41655 -15416 41768 -15380
rect 41721 -15434 41768 -15416
rect 73336 -15406 73713 -15372
rect 73336 -15460 73718 -15406
rect 73798 -15426 73856 -15336
rect 73876 -15414 73878 -15348
rect 73336 -15511 73722 -15460
rect 73696 -15528 73722 -15511
rect 73798 -15528 73856 -15494
rect 73975 -15528 73990 -15234
rect 73997 -15528 74044 -15180
rect 74009 -15562 74024 -15528
rect 74446 -15593 74481 -15587
rect 74759 -15675 74794 -15641
rect 74760 -15694 74794 -15675
rect 74779 -15935 74794 -15694
rect 74813 -15728 74848 -15694
rect 74813 -15935 74847 -15728
rect 74813 -15969 74828 -15935
<< metal1 >>
rect -2400 3800 -2200 4000
rect -2400 3400 -2200 3600
rect -2400 3000 -2200 3200
rect -2400 2600 -2200 2800
rect -2400 2200 -2200 2400
rect -2400 1800 -2200 2000
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XDD1
timestamp 1722639531
transform 1 0 73843 0 1 -15381
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XDD2
timestamp 1722639531
transform 1 0 74647 0 1 -15788
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XDD3
timestamp 1722639531
transform 1 0 74960 0 1 -15841
box -183 -183 183 183
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM1
timestamp 1722639531
transform 1 0 38150 0 1 -13741
box -903 -647 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM2
timestamp 1722639531
transform 1 0 38641 0 1 -14095
box -903 -647 278 358
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM3
timestamp 1722639531
transform 1 0 39211 0 1 -14440
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM4
timestamp 1722639531
transform 1 0 -20221 0 1 -11198
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM5
timestamp 1722639531
transform 1 0 -19542 0 1 -11293
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM6
timestamp 1722639531
transform 1 0 39890 0 1 -14535
box -387 -397 387 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM7
timestamp 1722639531
transform 1 0 40490 0 1 -14639
box -903 -647 278 358
use sky130_fd_pr__nfet_03v3_nvt_UNEQ2N  XM8
timestamp 1722639531
transform 1 0 40981 0 1 -14993
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM9
timestamp 1722639531
transform 1 0 -18942 0 1 -11397
box -903 -647 278 358
use sky130_fd_pr__nfet_g5v0d10v5_H7BQ24  XM10
timestamp 1722639531
transform 1 0 -18214 0 1 -11751
box -941 -628 515 358
use sky130_fd_pr__nfet_03v3_nvt_UNEQ2N  XM11
timestamp 1722639531
transform 1 0 41472 0 1 -15058
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_54RBUL  XM12
timestamp 1722639531
transform 1 0 57684 0 1 -15114
box -16029 -397 16029 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM13
timestamp 1722639531
transform 1 0 74239 0 1 -15271
box -903 -647 278 358
use sky130_fd_pr__pfet_g5v0d10v5_54RBUL  XM20
timestamp 1722639531
transform 1 0 -1416 0 1 -12130
box -16029 -397 16029 397
use sky130_fd_pr__nfet_g5v0d10v5_A3MY9Q  XM22
timestamp 1722639531
transform 1 0 24227 0 1 -12234
box -9679 -358 9679 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM24
timestamp 1722639531
transform 1 0 34119 0 1 -12299
box -903 -647 278 358
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM25
timestamp 1722639531
transform 1 0 34610 0 1 -12644
box -308 -397 308 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM26
timestamp 1722639531
transform 1 0 35210 0 1 -12739
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM27
timestamp 1722639531
transform 1 0 35889 0 1 -12834
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM28
timestamp 1722639531
transform 1 0 36568 0 1 -12929
box -387 -397 387 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM29
timestamp 1722639531
transform 1 0 37168 0 1 -13033
box -903 -647 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM30
timestamp 1722639531
transform 1 0 37659 0 1 -13387
box -903 -647 278 358
use sky130_fd_pr__res_xhigh_po_0p35_E5287M  XR1
timestamp 1722639531
transform 1 0 -17551 0 1 -1850
box -201 -10582 201 10582
use sky130_fd_pr__res_xhigh_po_0p35_7R768E  XR2
timestamp 0
transform 1 0 75291 0 1 -15445
box -201 -632 201 632
<< labels >>
flabel metal1 -2400 3800 -2200 4000 0 FreeSans 25600 0 0 0 vdd
port 0 nsew
flabel metal1 -2400 3400 -2200 3600 0 FreeSans 25600 0 0 0 vss
port 1 nsew
flabel metal1 -2400 3000 -2200 3200 0 FreeSans 25600 0 0 0 out
port 2 nsew
flabel metal1 -2400 2600 -2200 2800 0 FreeSans 25600 0 0 0 inm
port 3 nsew
flabel metal1 -2400 2200 -2200 2400 0 FreeSans 25600 0 0 0 inp
port 4 nsew
flabel metal1 -2400 1800 -2200 2000 0 FreeSans 25600 0 0 0 ena
port 5 nsew
<< end >>
