magic
tech sky130A
magscale 1 2
timestamp 1723585349
<< pwell >>
rect -201 -683 201 683
<< psubdiff >>
rect -165 613 -69 647
rect 69 613 165 647
rect -165 551 -131 613
rect 131 551 165 613
rect -165 -613 -131 -551
rect 131 -613 165 -551
rect -165 -647 -69 -613
rect 69 -647 165 -613
<< psubdiffcont >>
rect -69 613 69 647
rect -165 -551 -131 551
rect 131 -551 165 551
rect -69 -647 69 -613
<< xpolycontact >>
rect -35 85 35 517
rect -35 -517 35 -85
<< xpolyres >>
rect -35 -85 35 85
<< locali >>
rect -165 613 -69 647
rect 69 613 165 647
rect -165 551 -131 613
rect 131 551 165 613
rect -165 -613 -131 -551
rect 131 -613 165 -551
rect -165 -647 -69 -613
rect 69 -647 165 -613
<< viali >>
rect -19 102 19 499
rect -19 -499 19 -102
<< metal1 >>
rect -25 499 25 511
rect -25 102 -19 499
rect 19 102 25 499
rect -25 90 25 102
rect -25 -102 25 -90
rect -25 -499 -19 -102
rect 19 -499 25 -102
rect -25 -511 25 -499
<< properties >>
string FIXED_BBOX -148 -630 148 630
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.013 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 2.402k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
