magic
tech sky130A
magscale 1 2
timestamp 1723501348
<< locali >>
rect 11242 16406 11550 16408
rect -21003 16400 11550 16406
rect -21003 16397 11481 16400
rect 11534 16397 11550 16400
rect -21003 16384 -20989 16397
rect -21003 16229 -20990 16384
rect 11535 16348 11550 16397
rect -29810 15696 -27543 15700
rect -24220 15698 -22598 15700
rect -21001 15698 -20990 16229
rect -26973 15696 -22598 15698
rect -22440 15696 -20990 15698
rect -29810 15674 -20990 15696
rect -20926 16229 11481 16348
rect -29810 15673 -21023 15674
rect -29810 15672 -22640 15673
rect -29810 15562 -29542 15672
rect -20926 15662 -20588 16229
rect 11242 15662 11481 16229
rect -29810 15560 -24237 15562
rect -29810 15558 -22640 15560
rect -29810 15555 -21052 15558
rect -20926 15555 11481 15662
rect -29810 15373 11481 15555
rect -29810 15365 -26601 15373
rect -29810 14604 -27541 15365
rect -28028 14602 -27541 14604
rect -27150 14601 -26601 15365
rect -26056 15371 -25550 15373
rect -24421 15371 11481 15373
rect -26056 14801 -25555 15371
rect -26057 14762 -25555 14801
rect -26056 14579 -25555 14762
rect -24421 14579 -23938 15371
rect -26056 14578 -25585 14579
rect -24220 14578 -23938 14579
rect -22806 15368 11481 15371
rect -26056 14575 -26020 14578
rect -22806 14576 -22323 15368
rect -22621 14572 -22323 14576
rect -21188 15124 11481 15368
rect -21188 14636 -20588 15124
rect -21188 14573 -20584 14636
rect -21188 14572 -20988 14573
rect -20776 14554 -20584 14573
rect 11228 14554 11481 15124
rect -20776 14425 11481 14554
rect -20776 14424 11112 14425
rect 11229 14424 11481 14425
rect 11534 15497 11550 16348
rect 11534 15251 11546 15497
rect -20776 14386 -20545 14424
rect 11534 14393 11547 15251
rect 11532 14386 11547 14393
rect -20776 14385 11112 14386
rect 11229 14385 11547 14386
rect -20776 14357 11547 14385
rect -29806 14339 -29627 14342
rect -29806 14239 -27004 14339
rect -29806 13973 -29627 14239
rect -29806 13934 -27006 13973
rect -8615 13942 -8279 14357
rect -29806 13738 -29669 13934
rect -8610 13896 -8279 13942
rect -22987 13744 -22818 13745
rect -25810 13741 -25750 13743
rect -29806 13711 -26954 13738
rect -29803 13690 -26954 13711
rect -29803 13355 -29157 13690
rect -29800 13144 -29674 13355
rect -29455 13144 -29162 13355
rect -28782 13144 -28450 13690
rect -27167 13144 -26954 13690
rect -29800 13142 -26954 13144
rect -26562 13142 -26365 13740
rect -25973 13142 -25750 13741
rect -29800 13128 -25750 13142
rect -24935 13468 -24716 13744
rect -24490 13468 -24302 13744
rect -24078 13468 -23844 13744
rect -24935 13128 -23844 13468
rect -23026 13128 -22818 13744
rect -29800 13127 -22818 13128
rect -22001 13742 -21851 13744
rect -22001 13127 -21713 13742
rect -29800 13112 -21713 13127
rect -2527 13112 -2316 13752
rect -29800 13008 -2316 13112
rect -29800 13006 -21872 13008
rect -29800 13002 -25842 13006
rect -29800 12913 -29545 13002
rect -26998 12917 -25842 12918
rect -24799 12917 -23972 12918
rect -22949 12917 -21872 12918
rect -26998 12915 -21872 12917
rect -2342 12915 -2316 13008
rect -26998 12913 -2316 12915
rect -29800 12904 -2316 12913
rect -29800 12900 -26998 12904
rect -24806 12902 -2316 12904
rect -23947 12901 -2316 12902
rect -21854 12899 -2316 12901
rect -21851 12791 -21793 12899
rect -21851 12790 -21796 12791
<< viali >>
rect 11481 16397 11534 16400
rect -20989 16384 11535 16397
rect -20990 16348 11535 16384
rect -20990 15674 -20926 16348
rect -21023 15673 -20926 15674
rect -22640 15672 -20926 15673
rect -29542 15562 -20926 15672
rect -24237 15560 -20926 15562
rect -22640 15558 -20926 15560
rect -21052 15555 -20926 15558
rect 11112 14424 11229 14425
rect 11481 14424 11534 16348
rect -20545 14393 11534 14424
rect -20545 14386 11532 14393
rect 11112 14385 11229 14386
rect -21872 13006 -2342 13008
rect -25842 13002 -2342 13006
rect -29545 12918 -2342 13002
rect -29545 12913 -26998 12918
rect -25842 12917 -24799 12918
rect -23972 12917 -22949 12918
rect -21872 12915 -2342 12918
rect -23042 12793 -22987 12844
<< metal1 >>
rect 11475 16403 11540 16412
rect -21001 16400 11547 16403
rect -21001 16397 11481 16400
rect 11534 16397 11547 16400
rect -21001 16384 -20989 16397
rect -21001 16342 -20990 16384
rect 11535 16348 11547 16397
rect -20999 15692 -20990 16342
rect -22632 15691 -20990 15692
rect -24221 15690 -20990 15691
rect -26985 15689 -20990 15690
rect -29798 15674 -20990 15689
rect -20926 16334 11481 16348
rect -29798 15673 -21023 15674
rect -29798 15672 -22640 15673
rect -29798 15562 -29542 15672
rect -29798 15560 -24237 15562
rect -29798 15558 -22640 15560
rect -29798 15555 -21052 15558
rect -20926 15555 -20909 16334
rect -16462 16126 -16431 16127
rect -13303 16126 -13272 16127
rect -6662 16126 -6631 16127
rect -2871 16126 -2840 16127
rect -2714 16126 -2683 16127
rect -1766 16126 -1735 16127
rect -343 16126 -312 16127
rect 2342 16126 2373 16127
rect 3921 16126 3952 16127
rect 6291 16126 6322 16127
rect 8503 16126 8534 16127
rect -20429 16092 11081 16126
rect -20874 15796 -20806 15800
rect -20876 15744 -20866 15796
rect -20814 15744 -20804 15796
rect -29798 15546 -20909 15555
rect -29771 15464 -29571 15546
rect -27466 14948 -27429 15176
rect -27494 14896 -27484 14948
rect -27432 14896 -27422 14948
rect -27364 14905 -27331 15266
rect -27271 14998 -27235 15546
rect -26985 15541 -20909 15546
rect -26523 14993 -26488 15541
rect -24221 15540 -20909 15541
rect -26455 15226 -26445 15278
rect -26393 15226 -26383 15278
rect -26281 15226 -26271 15278
rect -26219 15226 -26209 15278
rect -26429 14942 -26394 15226
rect -27466 14404 -27429 14896
rect -26453 14890 -26443 14942
rect -26391 14890 -26381 14942
rect -26269 14941 -26234 15226
rect -25396 15218 -25386 15270
rect -25334 15218 -25324 15270
rect -25237 15220 -25227 15272
rect -25175 15220 -25165 15272
rect -24810 15222 -24800 15274
rect -24748 15222 -24738 15274
rect -26428 14406 -26392 14890
rect -26284 14889 -26274 14941
rect -26222 14889 -26212 14941
rect -27484 14352 -27474 14404
rect -27422 14352 -27412 14404
rect -27297 14352 -27287 14404
rect -27235 14352 -27225 14404
rect -26447 14354 -26437 14406
rect -26385 14354 -26375 14406
rect -26272 14405 -26237 14889
rect -26176 14566 -26138 15170
rect -25482 14566 -25442 15172
rect -25374 14952 -25344 15218
rect -25216 14952 -25186 15220
rect -25396 14900 -25386 14952
rect -25334 14900 -25324 14952
rect -25239 14900 -25229 14952
rect -25177 14900 -25167 14952
rect -26186 14514 -26176 14566
rect -26124 14514 -26114 14566
rect -25502 14514 -25492 14566
rect -25440 14514 -25430 14566
rect -26292 14353 -26282 14405
rect -26230 14353 -26220 14405
rect -25393 14361 -25324 14900
rect -25122 14540 -25076 15174
rect -25122 14514 -25074 14540
rect -29535 13930 -29104 14138
rect -29545 13878 -29535 13930
rect -29104 13878 -29094 13930
rect -28912 13873 -28902 13925
rect -28850 13873 -28840 13925
rect -29095 13749 -29085 13801
rect -29033 13749 -29023 13801
rect -29598 13580 -29528 13582
rect -29602 13528 -29592 13580
rect -29540 13528 -29528 13580
rect -30146 13268 -29946 13357
rect -29598 13268 -29528 13528
rect -29083 13320 -29043 13749
rect -29006 13532 -28996 13584
rect -28944 13532 -28934 13584
rect -30146 13206 -29522 13268
rect -28987 13237 -28951 13532
rect -28892 13322 -28856 13873
rect -28400 13748 -28390 13800
rect -28338 13748 -28328 13800
rect -28379 13602 -28339 13748
rect -28403 13550 -28393 13602
rect -28341 13550 -28331 13602
rect -28379 13505 -28339 13550
rect -28295 13549 -28285 13601
rect -28233 13549 -28223 13601
rect -28137 13549 -28127 13601
rect -28075 13549 -28065 13601
rect -28379 13435 -28320 13505
rect -28335 13328 -28320 13435
rect -28277 13286 -28244 13549
rect -28293 13234 -28283 13286
rect -28231 13234 -28221 13286
rect -28117 13285 -28084 13549
rect -27976 13548 -27966 13600
rect -27914 13548 -27904 13600
rect -27817 13549 -27807 13601
rect -27755 13549 -27745 13601
rect -27956 13285 -27923 13548
rect -27799 13285 -27766 13549
rect -27396 13548 -27386 13600
rect -27334 13548 -27324 13600
rect -27721 13331 -27660 13506
rect -27481 13331 -27420 13506
rect -28136 13233 -28126 13285
rect -28074 13233 -28064 13285
rect -27976 13233 -27966 13285
rect -27914 13233 -27904 13285
rect -27818 13233 -27808 13285
rect -27756 13233 -27746 13285
rect -30146 13205 -29813 13206
rect -30146 13157 -29946 13205
rect -29598 13204 -29528 13206
rect -27707 13066 -27661 13331
rect -27481 13066 -27442 13331
rect -27375 13284 -27342 13548
rect -27279 13447 -27241 14352
rect -25407 14309 -25397 14361
rect -25319 14309 -25309 14361
rect -26091 13932 -26055 13936
rect -26801 13849 -26791 13901
rect -26739 13849 -26729 13901
rect -26776 13800 -26742 13849
rect -26207 13843 -26197 13895
rect -26145 13843 -26135 13895
rect -26100 13880 -26090 13932
rect -26038 13880 -26028 13932
rect -25120 13898 -25074 14514
rect -26677 13803 -26645 13809
rect -26804 13748 -26794 13800
rect -26742 13748 -26732 13800
rect -26696 13751 -26686 13803
rect -26634 13751 -26624 13803
rect -27393 13232 -27383 13284
rect -27331 13232 -27321 13284
rect -26878 13072 -26838 13506
rect -26776 13246 -26742 13748
rect -26677 13328 -26645 13751
rect -26183 13686 -26154 13843
rect -26290 13072 -26250 13505
rect -26183 13246 -26153 13686
rect -26091 13330 -26055 13880
rect -25694 13840 -25684 13892
rect -25632 13840 -25622 13892
rect -25136 13846 -25126 13898
rect -25074 13846 -25064 13898
rect -24900 13859 -24854 15174
rect -24788 14947 -24758 15222
rect -24651 15217 -24641 15269
rect -24589 15217 -24579 15269
rect -23780 15220 -23770 15272
rect -23718 15220 -23708 15272
rect -23622 15222 -23612 15274
rect -23560 15222 -23550 15274
rect -24634 14948 -24604 15217
rect -24811 14938 -24801 14947
rect -24814 14895 -24801 14938
rect -24749 14895 -24739 14947
rect -24653 14896 -24643 14948
rect -24591 14896 -24581 14948
rect -24814 14450 -24739 14895
rect -24534 14564 -24494 15170
rect -23862 14939 -23826 15172
rect -23761 14948 -23727 15220
rect -23780 14939 -23770 14948
rect -23862 14905 -23770 14939
rect -23862 14620 -23826 14905
rect -23780 14896 -23770 14905
rect -23718 14896 -23708 14948
rect -23602 14947 -23568 15222
rect -23504 14997 -23471 15540
rect -23276 14997 -23243 15540
rect -22632 15537 -20909 15540
rect -23196 15222 -23186 15274
rect -23134 15222 -23124 15274
rect -23039 15222 -23029 15274
rect -22977 15222 -22967 15274
rect -22163 15224 -22153 15276
rect -22101 15224 -22091 15276
rect -22006 15228 -21996 15280
rect -21944 15228 -21934 15280
rect -23175 14949 -23141 15222
rect -23018 14949 -22984 15222
rect -23621 14895 -23611 14947
rect -23559 14895 -23549 14947
rect -23196 14897 -23186 14949
rect -23134 14897 -23124 14949
rect -23037 14897 -23027 14949
rect -22975 14897 -22965 14949
rect -22922 14686 -22886 15175
rect -22253 14936 -22205 15172
rect -22143 14953 -22111 15224
rect -21985 14954 -21953 15228
rect -21890 14994 -21860 15537
rect -21654 14992 -21624 15537
rect -20999 15535 -20909 15537
rect -21056 15338 -21046 15390
rect -20994 15338 -20984 15390
rect -21574 15219 -21564 15271
rect -21512 15219 -21502 15271
rect -21420 15219 -21410 15271
rect -21358 15219 -21348 15271
rect -22161 14936 -22151 14953
rect -22253 14903 -22151 14936
rect -22941 14634 -22931 14686
rect -22879 14634 -22869 14686
rect -23874 14568 -23864 14620
rect -23812 14568 -23802 14620
rect -23602 14570 -23592 14622
rect -23540 14570 -23530 14622
rect -22922 14586 -22886 14634
rect -24556 14512 -24546 14564
rect -24494 14512 -24484 14564
rect -23862 14562 -23826 14568
rect -24824 14398 -24814 14450
rect -24736 14398 -24726 14450
rect -24237 14396 -24227 14448
rect -24149 14396 -24139 14448
rect -24652 14302 -24642 14354
rect -24564 14302 -24554 14354
rect -25672 13586 -25636 13840
rect -25052 13768 -25042 13820
rect -24990 13768 -24980 13820
rect -24916 13768 -24906 13859
rect -24854 13768 -24844 13859
rect -25702 13534 -25692 13586
rect -25640 13534 -25630 13586
rect -25580 13540 -25570 13592
rect -25518 13540 -25508 13592
rect -25174 13542 -25164 13594
rect -25112 13542 -25102 13594
rect -25672 13314 -25636 13534
rect -25574 13278 -25538 13540
rect -25590 13226 -25580 13278
rect -25528 13226 -25518 13278
rect -27052 13071 -25754 13072
rect -25470 13071 -25436 13492
rect -25244 13071 -25210 13492
rect -25148 13276 -25112 13542
rect -25046 13316 -25000 13768
rect -24639 13613 -24567 14302
rect -24637 13551 -24569 13613
rect -24225 13605 -24152 14396
rect -23782 13758 -23772 13810
rect -23720 13758 -23710 13810
rect -24225 13549 -24154 13605
rect -23764 13314 -23728 13758
rect -25164 13224 -25154 13276
rect -25102 13224 -25092 13276
rect -23665 13270 -23633 13574
rect -23568 13317 -23538 14570
rect -23347 14534 -23337 14586
rect -23285 14534 -23275 14586
rect -22942 14534 -22932 14586
rect -22880 14534 -22870 14586
rect -22253 14563 -22205 14903
rect -22161 14901 -22151 14903
rect -22099 14901 -22089 14953
rect -22003 14902 -21993 14954
rect -21941 14902 -21931 14954
rect -21560 14945 -21528 15219
rect -21579 14893 -21569 14945
rect -21517 14893 -21507 14945
rect -21401 14943 -21369 15219
rect -21421 14891 -21411 14943
rect -21359 14891 -21349 14943
rect -21308 14578 -21260 15171
rect -23332 13298 -23302 14534
rect -22922 14528 -22886 14534
rect -22559 14505 -22549 14557
rect -22497 14505 -22487 14557
rect -22271 14511 -22261 14563
rect -22209 14511 -22199 14563
rect -22651 14348 -22587 14350
rect -22655 14296 -22645 14348
rect -22593 14296 -22583 14348
rect -22760 13878 -22750 13930
rect -22698 13878 -22688 13930
rect -23146 13806 -23110 13808
rect -23164 13754 -23154 13806
rect -23102 13754 -23092 13806
rect -23687 13218 -23677 13270
rect -23625 13218 -23615 13270
rect -23240 13269 -23208 13575
rect -23146 13314 -23110 13754
rect -22744 13315 -22705 13878
rect -22651 13541 -22587 14296
rect -23261 13217 -23251 13269
rect -23199 13217 -23189 13269
rect -22639 13231 -22611 13541
rect -22544 13315 -22502 14505
rect -22213 14479 -22121 14481
rect -22213 14470 -22150 14479
rect -22214 14426 -22150 14470
rect -22098 14426 -22088 14479
rect -21308 14465 -21259 14578
rect -22214 14425 -22112 14426
rect -22331 14331 -22321 14383
rect -22269 14331 -22259 14383
rect -22317 13313 -22275 14331
rect -22214 13540 -22171 14425
rect -21309 14389 -21259 14465
rect -21320 14337 -21310 14389
rect -21258 14337 -21248 14389
rect -21050 14386 -20998 15338
rect -20874 14633 -20806 15744
rect -20512 15524 -20472 16034
rect -20412 15808 -20381 16092
rect -20432 15756 -20422 15808
rect -20370 15798 -20360 15808
rect -20252 15798 -20221 16092
rect -20093 15798 -20062 16092
rect -19940 15798 -19909 16092
rect -19779 15798 -19748 16092
rect -19620 15798 -19589 16092
rect -19463 15798 -19432 16092
rect -19305 15798 -19274 16092
rect -19148 15798 -19117 16092
rect -18988 15798 -18957 16092
rect -18831 15798 -18800 16092
rect -18672 15798 -18641 16092
rect -18515 15798 -18484 16092
rect -18355 15798 -18324 16092
rect -18196 15798 -18165 16092
rect -18043 15798 -18012 16092
rect -17881 15798 -17850 16092
rect -17724 15798 -17693 16092
rect -17566 15798 -17535 16092
rect -17409 15798 -17378 16092
rect -17249 15798 -17218 16092
rect -17093 15798 -17062 16092
rect -16934 15798 -16903 16092
rect -16776 15798 -16745 16092
rect -16621 15798 -16590 16092
rect -16462 15798 -16431 16092
rect -16305 15798 -16274 16092
rect -16144 15798 -16113 16092
rect -15987 15798 -15956 16092
rect -15829 15798 -15798 16092
rect -15672 15798 -15641 16092
rect -15514 15798 -15483 16092
rect -15358 15798 -15327 16092
rect -15196 15798 -15165 16092
rect -15039 15798 -15008 16092
rect -14880 15798 -14849 16092
rect -14721 15798 -14690 16092
rect -14564 15798 -14533 16092
rect -14406 15798 -14375 16092
rect -14250 15798 -14219 16092
rect -14091 15798 -14060 16092
rect -13933 15798 -13902 16092
rect -13775 15798 -13744 16092
rect -13618 15798 -13587 16092
rect -13459 15798 -13428 16092
rect -13303 15798 -13272 16092
rect -13142 15798 -13111 16092
rect -12984 15798 -12953 16092
rect -12826 15798 -12795 16092
rect -12668 15798 -12637 16092
rect -12509 15798 -12478 16092
rect -12351 15798 -12320 16092
rect -12193 15798 -12162 16092
rect -12036 15798 -12005 16092
rect -11878 15798 -11847 16092
rect -11720 15798 -11689 16092
rect -11562 15798 -11531 16092
rect -11405 15798 -11374 16092
rect -11245 15798 -11214 16092
rect -11086 15798 -11055 16092
rect -10931 15798 -10900 16092
rect -10772 15798 -10741 16092
rect -10616 15798 -10585 16092
rect -10456 15798 -10425 16092
rect -10301 15798 -10270 16092
rect -10141 15798 -10110 16092
rect -9983 15798 -9952 16092
rect -9823 15798 -9792 16092
rect -9670 15798 -9639 16092
rect -9509 15798 -9478 16092
rect -9350 15798 -9319 16092
rect -9195 15798 -9164 16092
rect -9034 15798 -9003 16092
rect -8876 15798 -8845 16092
rect -8719 15798 -8688 16092
rect -8563 15798 -8532 16092
rect -8403 15798 -8372 16092
rect -8246 15798 -8215 16092
rect -8087 15798 -8056 16092
rect -7928 15798 -7897 16092
rect -7770 15798 -7739 16092
rect -7612 15798 -7581 16092
rect -7454 15798 -7423 16092
rect -7295 15798 -7264 16092
rect -7139 15798 -7108 16092
rect -6979 15798 -6948 16092
rect -6822 15798 -6791 16092
rect -6662 15798 -6631 16092
rect -6505 15798 -6474 16092
rect -6349 15798 -6318 16092
rect -6189 15798 -6158 16092
rect -6032 15798 -6001 16092
rect -5873 15798 -5842 16092
rect -5715 15798 -5684 16092
rect -5556 15798 -5525 16092
rect -5401 15798 -5370 16092
rect -5241 15798 -5210 16092
rect -5085 15798 -5054 16092
rect -4925 15798 -4894 16092
rect -4769 15798 -4738 16092
rect -4612 15798 -4581 16092
rect -4454 15798 -4423 16092
rect -4292 15798 -4261 16092
rect -4136 15798 -4105 16092
rect -3977 15798 -3946 16092
rect -3822 15798 -3791 16092
rect -3662 15798 -3631 16092
rect -3504 15798 -3473 16092
rect -3348 15798 -3317 16092
rect -3188 15798 -3157 16092
rect -3030 15798 -2999 16092
rect -2871 15798 -2840 16092
rect -2714 15798 -2683 16092
rect -2558 15798 -2527 16092
rect -2400 15798 -2369 16092
rect -2240 15798 -2209 16092
rect -2085 15798 -2054 16092
rect -1924 15798 -1893 16092
rect -1766 15798 -1735 16092
rect -1607 15798 -1576 16092
rect -1451 15798 -1420 16092
rect -1293 15798 -1262 16092
rect -1134 15798 -1103 16092
rect -974 15798 -943 16092
rect -818 15798 -787 16092
rect -660 15798 -629 16092
rect -505 15798 -474 16092
rect -343 15798 -312 16092
rect -185 15798 -154 16092
rect -29 15798 2 16092
rect 129 15798 160 16092
rect 288 15798 319 16092
rect 446 15798 477 16092
rect 605 15798 636 16092
rect 762 15798 793 16092
rect 921 15798 952 16092
rect 1078 15798 1109 16092
rect 1235 15798 1266 16092
rect 1392 15798 1423 16092
rect 1553 15798 1584 16092
rect 1708 15798 1739 16092
rect 1869 15798 1900 16092
rect 2027 15798 2058 16092
rect 2181 15798 2212 16092
rect 2342 15798 2373 16092
rect 2501 15798 2532 16092
rect 2659 15798 2690 16092
rect 2816 15798 2847 16092
rect 2973 15798 3004 16092
rect 3132 15798 3163 16092
rect 3290 15798 3321 16092
rect 3447 15798 3478 16092
rect 3607 15798 3638 16092
rect 3764 15798 3795 16092
rect 3921 15798 3952 16092
rect 4078 15798 4109 16092
rect 4237 15798 4268 16092
rect 4395 15798 4426 16092
rect 4553 15798 4584 16092
rect 4711 15798 4742 16092
rect 4868 15798 4899 16092
rect 5028 15798 5059 16092
rect 5187 15798 5218 16092
rect 5341 15798 5372 16092
rect 5502 15798 5533 16092
rect 5660 15798 5691 16092
rect 5818 15798 5849 16092
rect 5977 15798 6008 16092
rect 6134 15798 6165 16092
rect 6291 15798 6322 16092
rect 6450 15798 6481 16092
rect 6609 15798 6640 16092
rect 6766 15798 6797 16092
rect 6924 15798 6955 16092
rect 7083 15798 7114 16092
rect 7240 15798 7271 16092
rect 7397 15798 7428 16092
rect 7557 15798 7588 16092
rect 7714 15798 7745 16092
rect 7874 15798 7905 16092
rect 8031 15798 8062 16092
rect 8188 15798 8219 16092
rect 8346 15798 8377 16092
rect 8503 15798 8534 16092
rect 8662 15798 8693 16092
rect 8821 15798 8852 16092
rect 8978 15798 9009 16092
rect 9136 15798 9167 16092
rect 9293 15798 9324 16092
rect 9450 15798 9481 16092
rect 9610 15798 9641 16092
rect 9769 15798 9800 16092
rect 9926 15798 9957 16092
rect 10084 15798 10115 16092
rect 10241 15798 10272 16092
rect 10401 15798 10432 16092
rect 10557 15798 10588 16092
rect 10714 15798 10745 16092
rect 10873 15798 10904 16092
rect 11031 15798 11062 16092
rect 11125 15846 11158 16334
rect -20370 15764 11080 15798
rect -20370 15756 -20360 15764
rect -19620 15763 -19589 15764
rect -15196 15763 -15165 15764
rect -9983 15763 -9952 15764
rect -20525 15472 -20515 15524
rect -20463 15472 -20453 15524
rect 11080 15472 11090 15524
rect 11142 15472 11152 15524
rect -20426 15385 -20391 15396
rect -20445 15333 -20435 15385
rect -20383 15333 -20373 15385
rect -20426 15034 -20391 15333
rect 11112 15120 11141 15472
rect -20447 14982 -20437 15034
rect -20385 15019 -20375 15034
rect -20285 15019 11067 15020
rect -20385 14986 11067 15019
rect -20385 14985 -20217 14986
rect -20385 14982 -20375 14985
rect -20525 14431 -20489 14926
rect -20425 14692 -20392 14982
rect -20267 14692 -20234 14985
rect -20109 14692 -20076 14986
rect -19952 14692 -19919 14986
rect -19792 14692 -19759 14986
rect -19635 14692 -19602 14986
rect -19475 14692 -19442 14986
rect -19319 14692 -19286 14986
rect -19160 14692 -19127 14986
rect -19003 14692 -18970 14986
rect -18844 14692 -18811 14986
rect -18686 14692 -18653 14986
rect -18528 14692 -18495 14986
rect -18372 14692 -18339 14986
rect -18212 14692 -18179 14986
rect -18056 14692 -18023 14986
rect -17897 14692 -17864 14986
rect -17739 14692 -17706 14986
rect -17583 14692 -17550 14986
rect -17424 14692 -17391 14986
rect -17264 14692 -17231 14986
rect -17106 14692 -17073 14986
rect -16947 14692 -16914 14986
rect -16790 14692 -16757 14986
rect -16634 14692 -16601 14986
rect -16473 14692 -16440 14986
rect -16316 14692 -16283 14986
rect -16160 14692 -16127 14986
rect -16003 14692 -15970 14986
rect -15843 14692 -15810 14986
rect -15686 14692 -15653 14986
rect -15528 14692 -15495 14986
rect -15368 14692 -15335 14986
rect -15210 14692 -15177 14986
rect -15054 14692 -15021 14986
rect -14896 14692 -14863 14986
rect -14738 14692 -14705 14986
rect -14579 14692 -14546 14986
rect -14420 14692 -14387 14986
rect -14265 14692 -14232 14986
rect -14106 14692 -14073 14986
rect -13948 14692 -13915 14986
rect -13789 14692 -13756 14986
rect -13630 14692 -13597 14986
rect -13473 14692 -13440 14986
rect -13317 14692 -13284 14986
rect -13157 14692 -13124 14986
rect -12998 14692 -12965 14986
rect -12840 14692 -12807 14986
rect -12683 14692 -12650 14986
rect -12526 14692 -12493 14986
rect -12367 14692 -12334 14986
rect -12208 14692 -12175 14986
rect -12049 14692 -12016 14986
rect -11893 14692 -11860 14986
rect -11733 14692 -11700 14986
rect -11577 14692 -11544 14986
rect -11419 14692 -11386 14986
rect -11260 14692 -11227 14986
rect -11104 14692 -11071 14986
rect -10947 14692 -10914 14986
rect -10788 14692 -10755 14986
rect -10630 14692 -10597 14986
rect -10470 14692 -10437 14986
rect -10314 14692 -10281 14986
rect -10155 14692 -10122 14986
rect -9998 14692 -9965 14986
rect -9841 14692 -9808 14986
rect -9683 14692 -9650 14986
rect -9524 14692 -9491 14986
rect -9367 14692 -9334 14986
rect -9209 14692 -9176 14986
rect -9050 14692 -9017 14986
rect -8892 14692 -8859 14986
rect -8732 14692 -8699 14986
rect -8576 14692 -8543 14986
rect -8417 14692 -8384 14986
rect -8261 14692 -8228 14986
rect -8100 14692 -8067 14986
rect -7943 14692 -7910 14986
rect -7785 14692 -7752 14986
rect -7627 14692 -7594 14986
rect -7470 14692 -7437 14986
rect -7310 14692 -7277 14986
rect -7154 14692 -7121 14986
rect -6997 14692 -6964 14986
rect -6837 14692 -6804 14986
rect -6682 14692 -6649 14986
rect -6524 14692 -6491 14986
rect -6366 14692 -6333 14986
rect -6206 14692 -6173 14986
rect -6048 14692 -6015 14986
rect -5889 14692 -5856 14986
rect -5733 14692 -5700 14986
rect -5575 14692 -5542 14986
rect -5414 14692 -5381 14986
rect -5256 14692 -5223 14986
rect -5099 14692 -5066 14986
rect -4941 14692 -4908 14986
rect -4783 14692 -4750 14986
rect -4626 14692 -4593 14986
rect -4467 14692 -4434 14986
rect -4310 14692 -4277 14986
rect -4153 14692 -4120 14986
rect -3995 14692 -3962 14986
rect -3837 14692 -3804 14986
rect -3678 14692 -3645 14986
rect -3520 14692 -3487 14986
rect -3362 14692 -3329 14986
rect -3202 14692 -3169 14986
rect -3048 14692 -3015 14986
rect -2887 14692 -2854 14986
rect -2730 14692 -2697 14986
rect -2573 14692 -2540 14986
rect -2414 14692 -2381 14986
rect -2256 14692 -2223 14986
rect -2098 14692 -2065 14986
rect -1939 14692 -1906 14986
rect -1783 14692 -1750 14986
rect -1627 14692 -1594 14986
rect -1466 14692 -1433 14986
rect -1308 14692 -1275 14986
rect -1150 14692 -1117 14986
rect -991 14692 -958 14986
rect -833 14692 -800 14986
rect -676 14692 -643 14986
rect -517 14692 -484 14986
rect -359 14692 -326 14986
rect -201 14692 -168 14986
rect -44 14692 -11 14986
rect 114 14692 147 14986
rect 274 14692 307 14986
rect 430 14692 463 14986
rect 588 14692 621 14986
rect 746 14692 779 14986
rect 904 14692 937 14986
rect 1063 14692 1096 14986
rect 1219 14692 1252 14986
rect 1376 14692 1409 14986
rect 1537 14692 1570 14986
rect 1694 14692 1727 14986
rect 1851 14692 1884 14986
rect 2010 14692 2043 14986
rect 2167 14692 2200 14986
rect 2326 14692 2359 14986
rect 2482 14692 2515 14986
rect 2643 14692 2676 14986
rect 2801 14692 2834 14986
rect 2958 14692 2991 14986
rect 3117 14692 3150 14986
rect 3275 14692 3308 14986
rect 3431 14692 3464 14986
rect 3591 14692 3624 14986
rect 3747 14692 3780 14986
rect 3907 14692 3940 14986
rect 4063 14692 4096 14986
rect 4222 14692 4255 14986
rect 4379 14692 4412 14986
rect 4537 14692 4570 14986
rect 4696 14692 4729 14986
rect 4853 14692 4886 14986
rect 5011 14692 5044 14986
rect 5170 14692 5203 14986
rect 5328 14692 5361 14986
rect 5487 14692 5520 14986
rect 5646 14692 5679 14986
rect 5802 14692 5835 14986
rect 5961 14692 5994 14986
rect 6117 14692 6150 14986
rect 6278 14692 6311 14986
rect 6436 14692 6469 14986
rect 6593 14692 6626 14986
rect 6752 14692 6785 14986
rect 6913 14692 6946 14986
rect 7065 14692 7098 14986
rect 7225 14692 7258 14986
rect 7384 14692 7417 14986
rect 7541 14692 7574 14986
rect 7698 14692 7731 14986
rect 7855 14692 7888 14986
rect 8016 14692 8049 14986
rect 8174 14692 8207 14986
rect 8331 14692 8364 14986
rect 8488 14692 8521 14986
rect 8645 14692 8678 14986
rect 8806 14692 8839 14986
rect 8962 14692 8995 14986
rect 9121 14692 9154 14986
rect 9277 14692 9310 14986
rect 9437 14692 9470 14986
rect 9596 14692 9629 14986
rect 9753 14692 9786 14986
rect 9911 14692 9944 14986
rect 10070 14692 10103 14986
rect 10227 14692 10260 14986
rect 10384 14692 10417 14986
rect 10543 14692 10576 14986
rect 10698 14692 10731 14986
rect 10856 14692 10889 14986
rect 11016 14692 11049 14986
rect 11112 14795 11146 15120
rect 11093 14743 11103 14795
rect 11155 14743 11165 14795
rect -20443 14658 11067 14692
rect -18528 14657 -18495 14658
rect -18056 14657 -18023 14658
rect -16316 14657 -16283 14658
rect -16003 14657 -15970 14658
rect -14265 14657 -14232 14658
rect -12367 14657 -12334 14658
rect -11733 14657 -11700 14658
rect -11419 14657 -11386 14658
rect -10155 14657 -10122 14658
rect -9998 14657 -9965 14658
rect -9209 14657 -9176 14658
rect -7627 14657 -7594 14658
rect -7310 14657 -7277 14658
rect -6997 14657 -6964 14658
rect -2414 14657 -2381 14658
rect -1308 14657 -1275 14658
rect -991 14657 -958 14658
rect 274 14657 307 14658
rect 588 14657 621 14658
rect 904 14657 937 14658
rect 1219 14657 1252 14658
rect 1376 14657 1409 14658
rect 3117 14657 3150 14658
rect 3907 14657 3940 14658
rect 4537 14657 4570 14658
rect 4853 14657 4886 14658
rect 5961 14657 5994 14658
rect 6752 14657 6785 14658
rect 7225 14657 7258 14658
rect 11456 14431 11481 16334
rect -20569 14425 11481 14431
rect -20569 14424 11112 14425
rect 11229 14424 11481 14425
rect 11534 16342 11547 16348
rect 11534 14430 11541 16342
rect -20569 14386 -20545 14424
rect 11534 14393 11544 14430
rect 11532 14386 11544 14393
rect -21065 14334 -21055 14386
rect -21003 14334 -20993 14386
rect -20569 14385 11112 14386
rect 11229 14385 11544 14386
rect -20569 14380 11544 14385
rect -20569 14376 11541 14380
rect -20569 14374 11113 14376
rect 11202 14374 11541 14376
rect -20569 14373 -20536 14374
rect -2654 14026 -2644 14078
rect -2592 14026 -2582 14078
rect -22140 13878 -22130 13930
rect -22078 13878 -22068 13930
rect -22211 13231 -22183 13540
rect -22117 13316 -22078 13878
rect -21559 13817 -21549 13869
rect -21497 13817 -21487 13869
rect -21539 13558 -21504 13817
rect -18696 13558 -18663 13559
rect -14427 13558 -14394 13559
rect -10796 13558 -10763 13559
rect -10003 13558 -9971 13559
rect -9846 13558 -9814 13559
rect -8582 13558 -8550 13559
rect -6684 13558 -6652 13559
rect -21556 13523 -2685 13558
rect -21634 13074 -21603 13475
rect -21539 13250 -21504 13523
rect -21538 13248 -21505 13250
rect -21376 13248 -21343 13523
rect -21223 13248 -21190 13523
rect -21063 13248 -21030 13523
rect -20905 13248 -20872 13523
rect -20747 13248 -20714 13523
rect -20587 13248 -20554 13523
rect -20432 13248 -20399 13523
rect -20274 13248 -20241 13523
rect -20114 13248 -20081 13523
rect -19958 13248 -19925 13523
rect -19799 13248 -19766 13523
rect -19643 13248 -19610 13523
rect -19485 13248 -19452 13523
rect -19325 13248 -19292 13523
rect -19166 13248 -19133 13523
rect -19008 13248 -18975 13523
rect -18852 13248 -18819 13523
rect -18696 13248 -18663 13523
rect -18536 13248 -18503 13523
rect -18378 13248 -18345 13523
rect -18219 13248 -18186 13523
rect -18061 13248 -18028 13523
rect -17904 13248 -17871 13523
rect -17746 13248 -17713 13523
rect -17588 13248 -17555 13523
rect -17428 13248 -17395 13523
rect -17272 13248 -17239 13523
rect -17113 13248 -17080 13523
rect -16955 13248 -16922 13523
rect -16798 13248 -16765 13523
rect -16639 13248 -16606 13523
rect -16482 13248 -16449 13523
rect -16324 13248 -16291 13523
rect -16167 13248 -16134 13523
rect -16010 13248 -15977 13523
rect -15848 13248 -15815 13523
rect -15693 13248 -15660 13523
rect -15534 13248 -15501 13523
rect -15377 13248 -15344 13523
rect -15219 13248 -15186 13523
rect -15060 13248 -15027 13523
rect -14901 13248 -14868 13523
rect -14744 13248 -14711 13523
rect -14585 13248 -14552 13523
rect -14427 13248 -14394 13523
rect -14271 13248 -14238 13523
rect -14111 13248 -14078 13523
rect -13954 13248 -13921 13523
rect -13795 13248 -13762 13523
rect -13637 13248 -13604 13523
rect -13481 13248 -13448 13523
rect -13322 13248 -13289 13523
rect -13163 13248 -13130 13523
rect -13006 13248 -12973 13523
rect -12847 13248 -12814 13523
rect -12690 13248 -12657 13523
rect -12531 13248 -12498 13523
rect -12374 13248 -12341 13523
rect -12215 13248 -12182 13523
rect -12059 13248 -12026 13523
rect -11901 13248 -11868 13523
rect -11744 13248 -11711 13523
rect -11585 13248 -11552 13523
rect -11425 13248 -11392 13523
rect -11266 13248 -11233 13523
rect -11109 13248 -11076 13523
rect -10953 13248 -10920 13523
rect -10796 13248 -10763 13523
rect -10639 13248 -10606 13523
rect -10477 13248 -10444 13523
rect -10321 13248 -10288 13523
rect -10161 13248 -10129 13523
rect -10003 13248 -9971 13523
rect -9846 13248 -9814 13523
rect -9687 13248 -9655 13523
rect -9530 13248 -9498 13523
rect -9371 13248 -9339 13523
rect -9213 13248 -9181 13523
rect -9055 13248 -9023 13523
rect -8897 13248 -8865 13523
rect -8739 13248 -8707 13523
rect -8582 13248 -8550 13523
rect -8423 13248 -8391 13523
rect -8266 13248 -8234 13523
rect -8108 13248 -8076 13523
rect -7950 13248 -7918 13523
rect -7790 13248 -7758 13523
rect -7634 13248 -7602 13523
rect -7475 13248 -7443 13523
rect -7315 13248 -7283 13523
rect -7159 13248 -7127 13523
rect -7000 13248 -6968 13523
rect -6844 13248 -6812 13523
rect -6684 13248 -6652 13523
rect -6526 13248 -6494 13523
rect -6369 13248 -6337 13523
rect -6211 13248 -6179 13523
rect -6053 13248 -6021 13523
rect -5895 13248 -5863 13523
rect -5739 13248 -5707 13523
rect -5578 13248 -5546 13523
rect -5421 13248 -5389 13523
rect -5262 13248 -5230 13523
rect -5103 13248 -5071 13523
rect -4945 13248 -4913 13523
rect -4787 13248 -4755 13523
rect -4630 13248 -4598 13523
rect -4473 13248 -4441 13523
rect -4316 13248 -4284 13523
rect -4155 13248 -4123 13523
rect -3999 13248 -3967 13523
rect -3841 13248 -3809 13523
rect -3682 13248 -3650 13523
rect -3527 13248 -3495 13523
rect -3366 13248 -3334 13523
rect -3208 13248 -3176 13523
rect -3051 13248 -3019 13523
rect -2892 13248 -2860 13523
rect -2736 13248 -2704 13523
rect -2641 13301 -2612 14026
rect -21554 13213 -2683 13248
rect -21857 13073 -2324 13074
rect -23957 13072 -2324 13073
rect -24802 13071 -2324 13072
rect -27052 13066 -2324 13071
rect -29801 13064 -28394 13066
rect -28335 13064 -2324 13066
rect -29801 13008 -2324 13064
rect -29801 13006 -21872 13008
rect -29801 13002 -25842 13006
rect -29801 12913 -29545 13002
rect -26998 12917 -25842 12918
rect -24799 12917 -23972 12918
rect -22949 12917 -21872 12918
rect -26998 12915 -21872 12917
rect -2342 12915 -2324 13008
rect -26998 12913 -2324 12915
rect -29801 12906 -2324 12913
rect -29801 12902 -21857 12906
rect -29801 12900 -25754 12902
rect -23957 12901 -21857 12902
rect -29801 12899 -26972 12900
rect -29771 12898 -29552 12899
rect -27008 12898 -26972 12899
rect -29771 12846 -29569 12898
rect -29771 12844 -29571 12846
rect -23059 12787 -23049 12850
rect -22978 12787 -22968 12850
<< via1 >>
rect -20866 15744 -20814 15796
rect -27484 14896 -27432 14948
rect -26445 15226 -26393 15278
rect -26271 15226 -26219 15278
rect -26443 14890 -26391 14942
rect -25386 15218 -25334 15270
rect -25227 15220 -25175 15272
rect -24800 15222 -24748 15274
rect -26274 14889 -26222 14941
rect -27474 14352 -27422 14404
rect -27287 14352 -27235 14404
rect -26437 14354 -26385 14406
rect -25386 14900 -25334 14952
rect -25229 14900 -25177 14952
rect -26176 14514 -26124 14566
rect -25492 14514 -25440 14566
rect -26282 14353 -26230 14405
rect -29535 13878 -29104 13930
rect -28902 13873 -28850 13925
rect -29085 13749 -29033 13801
rect -29592 13528 -29540 13580
rect -28996 13532 -28944 13584
rect -28390 13748 -28338 13800
rect -28393 13550 -28341 13602
rect -28285 13549 -28233 13601
rect -28127 13549 -28075 13601
rect -28283 13234 -28231 13286
rect -27966 13548 -27914 13600
rect -27807 13549 -27755 13601
rect -27386 13548 -27334 13600
rect -28126 13233 -28074 13285
rect -27966 13233 -27914 13285
rect -27808 13233 -27756 13285
rect -25397 14309 -25319 14361
rect -26791 13849 -26739 13901
rect -26197 13843 -26145 13895
rect -26090 13880 -26038 13932
rect -26794 13748 -26742 13800
rect -26686 13751 -26634 13803
rect -27383 13232 -27331 13284
rect -25684 13840 -25632 13892
rect -25126 13846 -25074 13898
rect -24641 15217 -24589 15269
rect -23770 15220 -23718 15272
rect -23612 15222 -23560 15274
rect -24801 14895 -24749 14947
rect -24643 14896 -24591 14948
rect -23770 14896 -23718 14948
rect -23186 15222 -23134 15274
rect -23029 15222 -22977 15274
rect -22153 15224 -22101 15276
rect -21996 15228 -21944 15280
rect -23611 14895 -23559 14947
rect -23186 14897 -23134 14949
rect -23027 14897 -22975 14949
rect -21046 15338 -20994 15390
rect -21564 15219 -21512 15271
rect -21410 15219 -21358 15271
rect -22931 14634 -22879 14686
rect -23864 14568 -23812 14620
rect -23592 14570 -23540 14622
rect -24546 14512 -24494 14564
rect -24814 14398 -24736 14450
rect -24227 14396 -24149 14448
rect -24642 14302 -24564 14354
rect -25042 13768 -24990 13820
rect -24906 13768 -24854 13859
rect -25692 13534 -25640 13586
rect -25570 13540 -25518 13592
rect -25164 13542 -25112 13594
rect -25580 13226 -25528 13278
rect -23772 13758 -23720 13810
rect -25154 13224 -25102 13276
rect -23337 14534 -23285 14586
rect -22932 14534 -22880 14586
rect -22151 14901 -22099 14953
rect -21993 14902 -21941 14954
rect -21569 14893 -21517 14945
rect -21411 14891 -21359 14943
rect -22549 14505 -22497 14557
rect -22261 14511 -22209 14563
rect -22645 14296 -22593 14348
rect -22750 13878 -22698 13930
rect -23154 13754 -23102 13806
rect -23677 13218 -23625 13270
rect -23251 13217 -23199 13269
rect -22150 14426 -22098 14479
rect -22321 14331 -22269 14383
rect -21310 14337 -21258 14389
rect -20422 15756 -20370 15808
rect -20515 15472 -20463 15524
rect 11090 15472 11142 15524
rect -20435 15333 -20383 15385
rect -20437 14982 -20385 15034
rect 11103 14743 11155 14795
rect -21055 14334 -21003 14386
rect -2644 14026 -2592 14078
rect -22130 13878 -22078 13930
rect -21549 13817 -21497 13869
rect -23049 12844 -22978 12850
rect -23049 12793 -23042 12844
rect -23042 12793 -22987 12844
rect -22987 12793 -22978 12844
rect -23049 12787 -22978 12793
<< metal2 >>
rect -20422 15808 -20370 15818
rect -20866 15798 -20814 15806
rect -20874 15797 -20806 15798
rect -20874 15796 -20422 15797
rect -20874 15763 -20866 15796
rect -20814 15764 -20422 15796
rect -20814 15763 -20806 15764
rect -20370 15764 -20361 15797
rect -20422 15746 -20370 15756
rect -20866 15734 -20814 15744
rect -20515 15524 -20463 15534
rect 11090 15524 11142 15534
rect 11089 15517 11090 15521
rect -20463 15477 11090 15517
rect -20515 15462 -20463 15472
rect 11089 15472 11090 15477
rect 11598 15521 11806 15608
rect 11142 15472 11806 15521
rect 11089 15468 11806 15472
rect 11090 15462 11142 15468
rect -21046 15392 -20994 15400
rect 11598 15395 11806 15468
rect -20435 15392 -20383 15395
rect -21048 15390 -20375 15392
rect -21048 15338 -21046 15390
rect -20994 15385 -20375 15390
rect -20994 15338 -20435 15385
rect -21048 15334 -20435 15338
rect -21046 15328 -20994 15334
rect -20383 15334 -20375 15385
rect -20435 15323 -20383 15333
rect -26445 15278 -26393 15288
rect -26448 15228 -26445 15261
rect -26271 15278 -26219 15288
rect -26393 15228 -26271 15261
rect -26445 15216 -26393 15226
rect -25386 15270 -25334 15280
rect -25393 15233 -25386 15267
rect -26271 15216 -26219 15226
rect -25227 15272 -25175 15282
rect -25334 15233 -25227 15267
rect -25386 15208 -25334 15218
rect -24800 15274 -24748 15284
rect -25175 15233 -25165 15267
rect -24810 15233 -24800 15267
rect -25227 15210 -25175 15220
rect -24641 15269 -24589 15279
rect -24748 15233 -24641 15267
rect -24800 15212 -24748 15222
rect -23770 15272 -23718 15282
rect -24589 15233 -24582 15267
rect -23777 15234 -23770 15267
rect -24641 15207 -24589 15217
rect -23612 15274 -23560 15284
rect -23718 15234 -23612 15267
rect -23770 15210 -23718 15220
rect -23186 15274 -23134 15284
rect -23560 15234 -23186 15267
rect -23612 15212 -23560 15222
rect -23029 15274 -22977 15284
rect -23134 15234 -23029 15267
rect -23186 15212 -23134 15222
rect -22153 15276 -22101 15286
rect -22977 15234 -22967 15267
rect -22161 15228 -22153 15262
rect -23029 15212 -22977 15222
rect -21996 15280 -21944 15290
rect -22101 15228 -21996 15262
rect -21564 15271 -21512 15281
rect -21944 15228 -21564 15262
rect -22153 15214 -22101 15224
rect -21996 15218 -21944 15228
rect -21410 15271 -21358 15281
rect -21512 15228 -21410 15262
rect -21564 15209 -21512 15219
rect -21358 15228 -21349 15262
rect -21410 15209 -21358 15219
rect -20437 15034 -20385 15044
rect -20437 14972 -20385 14982
rect -27484 14948 -27432 14958
rect -25386 14952 -25334 14962
rect -26443 14942 -26391 14952
rect -27432 14904 -27314 14938
rect -26445 14903 -26443 14936
rect -27484 14886 -27432 14896
rect -26274 14941 -26222 14951
rect -26391 14903 -26274 14936
rect -26443 14880 -26391 14890
rect -26222 14903 -26220 14936
rect -25394 14906 -25386 14940
rect -25229 14952 -25177 14962
rect -25334 14906 -25229 14940
rect -25386 14890 -25334 14900
rect -24801 14947 -24749 14957
rect -25177 14906 -25166 14940
rect -24808 14906 -24801 14940
rect -25229 14890 -25177 14900
rect -24643 14948 -24591 14958
rect -24749 14906 -24643 14940
rect -26274 14879 -26222 14889
rect -24801 14885 -24749 14895
rect -23770 14948 -23718 14958
rect -24591 14906 -24580 14940
rect -23777 14906 -23770 14939
rect -24643 14886 -24591 14896
rect -23611 14947 -23559 14957
rect -23718 14906 -23611 14939
rect -23770 14886 -23718 14896
rect -23186 14949 -23134 14959
rect -23559 14906 -23186 14939
rect -23611 14885 -23559 14895
rect -23027 14949 -22975 14959
rect -23134 14906 -23027 14939
rect -23186 14887 -23134 14897
rect -22151 14953 -22099 14963
rect -22975 14906 -22967 14939
rect -22160 14903 -22151 14937
rect -23027 14887 -22975 14897
rect -21993 14954 -21941 14964
rect -22099 14903 -21993 14937
rect -22151 14891 -22099 14901
rect -21569 14945 -21517 14955
rect -21941 14903 -21569 14937
rect -21993 14892 -21941 14902
rect -21411 14943 -21359 14953
rect -21517 14903 -21411 14937
rect -21569 14883 -21517 14893
rect -21359 14903 -21348 14937
rect -21411 14881 -21359 14891
rect 11097 14805 11147 14821
rect 11097 14795 11155 14805
rect 11097 14743 11103 14795
rect 11097 14733 11155 14743
rect -22927 14696 -20807 14701
rect -22931 14686 -20807 14696
rect -22879 14635 -20807 14686
rect -23864 14625 -23812 14630
rect -23592 14625 -23540 14632
rect -23864 14622 -23537 14625
rect -22931 14624 -22879 14634
rect -23864 14620 -23592 14622
rect -26176 14566 -26124 14576
rect -25492 14566 -25440 14576
rect -24546 14566 -24494 14574
rect -26124 14514 -25492 14566
rect -25440 14564 -24494 14566
rect -25440 14514 -24546 14564
rect -26176 14504 -26124 14514
rect -25500 14512 -24546 14514
rect -23812 14570 -23592 14620
rect -23540 14570 -23537 14622
rect -23812 14568 -23537 14570
rect -23864 14562 -23537 14568
rect -23337 14590 -23285 14596
rect -22960 14590 -22880 14596
rect -23337 14586 -22880 14590
rect -23864 14558 -23812 14562
rect -23592 14560 -23540 14562
rect -23285 14534 -22932 14586
rect -23337 14524 -22880 14534
rect -22549 14557 -22497 14567
rect -22261 14563 -22209 14573
rect -25492 14504 -25440 14512
rect -24546 14502 -24494 14512
rect -22497 14512 -22261 14557
rect -22549 14495 -22497 14505
rect -22209 14512 -22205 14557
rect -22261 14501 -22209 14511
rect -22150 14479 -22098 14489
rect -24814 14450 -24736 14460
rect -24224 14458 -22150 14465
rect -27474 14404 -27422 14414
rect -27287 14404 -27235 14414
rect -27422 14365 -27287 14402
rect -27474 14342 -27422 14352
rect -26437 14406 -26385 14416
rect -27235 14364 -26437 14398
rect -27287 14342 -27235 14352
rect -26282 14405 -26230 14415
rect -24820 14405 -24814 14443
rect -26385 14364 -26282 14398
rect -26437 14344 -26385 14354
rect -24227 14448 -22150 14458
rect -24736 14405 -24227 14443
rect -24814 14388 -24736 14398
rect -24149 14428 -22150 14448
rect -22180 14427 -22150 14428
rect -22098 14427 -22093 14465
rect -22150 14416 -22098 14426
rect -24227 14386 -24149 14396
rect -22321 14385 -22269 14393
rect -21310 14390 -21258 14399
rect -21055 14390 -21003 14396
rect -21310 14389 -20998 14390
rect -22321 14383 -21310 14385
rect -26282 14343 -26230 14353
rect -25397 14361 -25319 14371
rect -24642 14354 -24564 14364
rect -25319 14312 -24642 14347
rect -25397 14299 -25319 14309
rect -22645 14349 -22593 14358
rect -24564 14348 -22588 14349
rect -24564 14302 -22645 14348
rect -24642 14296 -22645 14302
rect -22593 14296 -22588 14348
rect -22269 14337 -21310 14383
rect -21258 14386 -20998 14389
rect -21258 14337 -21055 14386
rect -22321 14321 -22269 14331
rect -21310 14335 -21055 14337
rect -21310 14327 -21258 14335
rect -21003 14335 -20998 14386
rect -21055 14324 -21003 14334
rect -24642 14294 -22588 14296
rect -24642 14292 -24564 14294
rect -22645 14286 -22593 14294
rect 11097 14090 11147 14733
rect 11094 14088 11147 14090
rect -2644 14078 11147 14088
rect -2592 14029 11147 14078
rect -2644 14016 -2592 14026
rect 11094 14018 11146 14029
rect -29535 13930 -29104 13940
rect -28902 13925 -28850 13935
rect -29104 13878 -28902 13921
rect -29535 13868 -29104 13878
rect -26090 13933 -26034 13943
rect -28902 13863 -28850 13873
rect -26791 13901 -26739 13911
rect -26197 13895 -26145 13905
rect -26739 13849 -26197 13892
rect -26791 13839 -26739 13849
rect -22753 13932 -22697 13942
rect -26090 13867 -26034 13877
rect -25684 13892 -25632 13902
rect -25126 13898 -25074 13908
rect -26197 13833 -26145 13843
rect -25632 13860 -25126 13892
rect -25684 13830 -25632 13840
rect -25126 13836 -25074 13846
rect -24906 13862 -24854 13869
rect -23830 13862 -23662 13878
rect -23212 13862 -23044 13874
rect -22753 13866 -22697 13876
rect -22132 13932 -22076 13942
rect -22132 13866 -22076 13876
rect -21549 13869 -21497 13879
rect -24906 13859 -22781 13862
rect -25042 13820 -24990 13830
rect -29085 13801 -29033 13811
rect -28390 13800 -28338 13810
rect -29033 13750 -28390 13800
rect -29085 13739 -29033 13749
rect -28396 13748 -28390 13750
rect -26794 13800 -26742 13810
rect -28338 13748 -26794 13796
rect -28390 13738 -28338 13748
rect -26794 13738 -26742 13748
rect -26688 13805 -26632 13815
rect -25046 13768 -25042 13806
rect -24990 13768 -24906 13806
rect -24854 13850 -22781 13859
rect -24854 13829 -23802 13850
rect -23690 13846 -22781 13850
rect -23690 13829 -23184 13846
rect -23072 13838 -22781 13846
rect -22669 13838 -22160 13862
rect -23072 13837 -22160 13838
rect -22047 13837 -21549 13862
rect -23072 13829 -21549 13837
rect -25042 13758 -24990 13768
rect -24906 13758 -24854 13768
rect -23774 13812 -23718 13822
rect -26688 13739 -26632 13749
rect -23774 13746 -23718 13756
rect -23156 13808 -23100 13818
rect -22809 13807 -22637 13829
rect -22195 13806 -22015 13829
rect -21549 13807 -21497 13817
rect -23156 13742 -23100 13752
rect -28393 13602 -28341 13612
rect -29592 13582 -29540 13590
rect -28996 13584 -28944 13594
rect -29600 13580 -28996 13582
rect -29600 13548 -29592 13580
rect -29540 13548 -28996 13580
rect -29592 13518 -29540 13528
rect -28944 13548 -28934 13582
rect -28285 13601 -28233 13611
rect -28292 13591 -28285 13594
rect -28341 13558 -28285 13591
rect -28393 13540 -28341 13550
rect -28127 13601 -28075 13611
rect -28233 13559 -28127 13594
rect -28285 13539 -28233 13549
rect -27966 13600 -27914 13610
rect -28075 13559 -27966 13594
rect -28127 13539 -28075 13549
rect -27807 13601 -27755 13611
rect -27914 13559 -27807 13594
rect -27966 13538 -27914 13548
rect -27386 13600 -27334 13610
rect -27755 13559 -27386 13594
rect -27807 13539 -27755 13549
rect -27334 13559 -27320 13594
rect -25692 13586 -25640 13596
rect -27386 13538 -27334 13548
rect -28996 13522 -28944 13532
rect -25570 13592 -25518 13602
rect -25640 13544 -25570 13578
rect -25588 13542 -25570 13544
rect -25692 13524 -25640 13534
rect -25164 13594 -25112 13604
rect -25518 13542 -25164 13576
rect -25112 13542 -25092 13576
rect -25570 13530 -25518 13540
rect -25164 13532 -25112 13542
rect -28283 13286 -28231 13296
rect -28290 13245 -28283 13280
rect -28126 13285 -28074 13295
rect -28231 13245 -28126 13280
rect -28283 13224 -28231 13234
rect -27966 13285 -27914 13295
rect -28074 13245 -27966 13280
rect -28126 13223 -28074 13233
rect -27808 13285 -27756 13295
rect -27914 13245 -27808 13280
rect -27966 13223 -27914 13233
rect -27383 13284 -27331 13294
rect -27756 13245 -27383 13280
rect -27808 13223 -27756 13233
rect -27331 13245 -27318 13280
rect -25580 13278 -25528 13288
rect -25588 13232 -25580 13266
rect -27383 13222 -27331 13232
rect -25154 13276 -25102 13286
rect -25528 13232 -25154 13266
rect -25580 13216 -25528 13226
rect -23677 13273 -23625 13280
rect -23251 13273 -23199 13279
rect -23698 13270 -23596 13273
rect -25102 13232 -25092 13266
rect -25154 13214 -25102 13224
rect -23698 13218 -23677 13270
rect -23625 13218 -23596 13270
rect -23698 12901 -23596 13218
rect -23272 13269 -23170 13273
rect -23272 13217 -23251 13269
rect -23199 13217 -23170 13269
rect -23272 12901 -23170 13217
rect -23699 12814 -23596 12901
rect -23273 12849 -23170 12901
rect -23049 12851 -22978 12860
rect -23079 12850 -22955 12851
rect -23079 12849 -23049 12850
rect -23273 12819 -23049 12849
rect -23751 12614 -23550 12814
rect -23335 12789 -23049 12819
rect -23335 12619 -23134 12789
rect -23079 12788 -23049 12789
rect -22978 12788 -22955 12850
rect -23049 12777 -22978 12787
<< via2 >>
rect -26090 13932 -26034 13933
rect -26090 13880 -26038 13932
rect -26038 13880 -26034 13932
rect -22753 13930 -22697 13932
rect -26090 13877 -26034 13880
rect -22753 13878 -22750 13930
rect -22750 13878 -22698 13930
rect -22698 13878 -22697 13930
rect -22753 13876 -22697 13878
rect -22132 13930 -22076 13932
rect -22132 13878 -22130 13930
rect -22130 13878 -22078 13930
rect -22078 13878 -22076 13930
rect -22132 13876 -22076 13878
rect -26688 13803 -26632 13805
rect -26688 13751 -26686 13803
rect -26686 13751 -26634 13803
rect -26634 13751 -26632 13803
rect -23774 13810 -23718 13812
rect -23774 13758 -23772 13810
rect -23772 13758 -23720 13810
rect -23720 13758 -23718 13810
rect -26688 13749 -26632 13751
rect -23774 13756 -23718 13758
rect -23156 13806 -23100 13808
rect -23156 13754 -23154 13806
rect -23154 13754 -23102 13806
rect -23102 13754 -23100 13806
rect -23156 13752 -23100 13754
<< metal3 >>
rect -26090 13940 -22098 13942
rect -26091 13938 -22098 13940
rect -26100 13937 -22098 13938
rect -26100 13933 -22066 13937
rect -26100 13877 -26090 13933
rect -26034 13932 -22066 13933
rect -26034 13880 -22753 13932
rect -26034 13877 -26024 13880
rect -26100 13872 -26024 13877
rect -22763 13876 -22753 13880
rect -22697 13880 -22132 13932
rect -22697 13876 -22687 13880
rect -22763 13871 -22687 13876
rect -22142 13876 -22132 13880
rect -22076 13876 -22066 13932
rect -22142 13871 -22066 13876
rect -23784 13812 -23708 13817
rect -26698 13808 -26622 13810
rect -23784 13808 -23774 13812
rect -26708 13805 -23774 13808
rect -26708 13749 -26688 13805
rect -26632 13756 -23774 13805
rect -23718 13808 -23708 13812
rect -23166 13808 -23090 13813
rect -23718 13756 -23156 13808
rect -26632 13752 -23156 13756
rect -23100 13752 -23090 13808
rect -26632 13749 -23090 13752
rect -26708 13748 -23090 13749
rect -26698 13744 -26622 13748
rect -23166 13747 -23090 13748
use sky130_fd_pr__res_generic_l1_DBPZV5  sky130_fd_pr__res_generic_l1_DBPZV5_0
timestamp 1723067318
transform 0 1 -22404 -1 0 12820
box -30 -610 30 610
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XDD1
timestamp 1723064828
transform 1 0 -24603 0 1 13581
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XDD2
timestamp 1723064828
transform 1 0 -29561 0 1 13240
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XDD3
timestamp 1723064828
transform 1 0 -24190 0 1 13581
box -183 -183 183 183
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM1
timestamp 1723064828
transform 1 0 -23648 0 1 13403
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM2
timestamp 1723064828
transform 1 0 -23222 0 1 13403
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM3
timestamp 1723064828
transform 1 0 -21464 0 1 15083
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM4
timestamp 1723064828
transform 1 0 -23080 0 1 15086
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM5
timestamp 1723064828
transform 1 0 -23664 0 1 15086
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM6
timestamp 1723064828
transform 1 0 -22048 0 1 15083
box -387 -397 387 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM7
timestamp 1723064828
transform 1 0 -26169 0 1 13417
box -278 -358 278 358
use sky130_fd_pr__nfet_03v3_nvt_UNEQ2N  XM8
timestamp 1723064828
transform 1 0 -22623 0 1 13403
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM9
timestamp 1723064828
transform 1 0 -26758 0 1 13417
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_H7BQ24  XM10
timestamp 1723064828
transform 1 0 -28020 0 1 13419
box -515 -358 515 358
use sky130_fd_pr__nfet_03v3_nvt_UNEQ2N  XM11
timestamp 1723064828
transform 1 0 -22197 0 1 13403
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_54RBUL  XM12
timestamp 1723064828
transform 1 0 -4674 0 1 15945
box -16029 -397 16029 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM13
timestamp 1723064828
transform 1 0 -28969 0 1 13409
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_54RBUL  XM20
timestamp 1723064828
transform 1 0 -4688 0 1 14839
box -16029 -397 16029 397
use sky130_fd_pr__nfet_g5v0d10v5_A3MY9Q  XM22
timestamp 1723064828
transform 1 0 -12120 0 1 13386
box -9679 -358 9679 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM24
timestamp 1723064828
transform 1 0 -27357 0 1 13419
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM25
timestamp 1723064828
transform 1 0 -27348 0 1 15085
box -308 -397 308 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM26
timestamp 1723064828
transform 1 0 -26332 0 1 15081
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM27
timestamp 1723064828
transform 1 0 -25280 0 1 15086
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM28
timestamp 1723064828
transform 1 0 -24696 0 1 15086
box -387 -397 387 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM29
timestamp 1723064828
transform 1 0 -25128 0 1 13405
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM30
timestamp 1723064828
transform 1 0 -25554 0 1 13405
box -278 -358 278 358
use sky130_fd_pr__res_xhigh_po_0p35_E5287M  XR1
timestamp 1723064828
transform 0 1 -19120 -1 0 14103
box -201 -10582 201 10582
use sky130_fd_pr__res_xhigh_po_0p35_7R768E  XR2
timestamp 0
transform 1 0 -22885 0 1 12615
box 0 0 1 1
<< labels >>
flabel metal1 -29771 12844 -29571 13044 0 FreeSans 480 0 0 0 vss
port 1 nsew
flabel metal2 -23749 12615 -23550 12814 0 FreeSans 480 0 0 0 inm
port 3 nsew
flabel metal2 -23334 12619 -23134 12818 0 FreeSans 480 0 0 0 inp
port 4 nsew
flabel metal1 -30146 13157 -29946 13357 0 FreeSans 480 0 0 0 ena
port 5 nsew
flabel metal1 -29771 15464 -29571 15664 0 FreeSans 480 0 0 0 vdd
port 0 nsew
flabel metal2 11602 15402 11802 15602 0 FreeSans 480 0 0 0 out
port 2 nsew
<< end >>
