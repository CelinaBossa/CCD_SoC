magic
tech sky130A
magscale 1 2
timestamp 1723587632
<< dnwell >>
rect -4467 -3821 2737 6561
<< nwell >>
rect -4547 6326 2817 6641
rect -4547 -3586 -4232 6326
rect 2502 -3586 2817 6326
rect -4547 -3901 2817 -3586
<< mvnsubdiff >>
rect -4481 6555 2751 6575
rect -4481 6521 -4401 6555
rect 2671 6521 2751 6555
rect -4481 6501 2751 6521
rect -4481 6495 -4407 6501
rect -4481 -3755 -4461 6495
rect -4427 -3755 -4407 6495
rect -4481 -3761 -4407 -3755
rect 2677 6495 2751 6501
rect 2677 -3755 2697 6495
rect 2731 -3755 2751 6495
rect 2677 -3761 2751 -3755
rect -4481 -3781 2751 -3761
rect -4481 -3815 -4401 -3781
rect 2671 -3815 2751 -3781
rect -4481 -3835 2751 -3815
<< mvnsubdiffcont >>
rect -4401 6521 2671 6555
rect -4461 -3755 -4427 6495
rect 2697 -3755 2731 6495
rect -4401 -3815 2671 -3781
<< locali >>
rect -4461 6521 -4401 6555
rect 2671 6521 2731 6555
rect -4461 6495 2731 6521
rect -4462 -542 -4461 990
rect -4427 6488 2697 6495
rect -4427 6347 -4332 6488
rect 2644 6347 2697 6488
rect -4427 6298 2697 6347
rect -4427 4172 -4344 6298
rect -4257 6252 2697 6298
rect -4257 4172 -4147 6252
rect -4427 3929 -4147 4172
rect 2432 3929 2697 6252
rect -4427 3889 -4150 3929
rect 2440 3889 2697 3929
rect -4427 1567 -4147 3889
rect 2432 1567 2697 3889
rect -4427 1432 2697 1567
rect -4427 1431 2127 1432
rect -4427 1190 -4064 1431
rect -3828 1410 2127 1431
rect -3828 1190 -3415 1410
rect -4427 1182 -3415 1190
rect -4427 1120 -4349 1182
rect -4156 1177 -3415 1182
rect -4156 1120 -4140 1177
rect -4427 164 -4140 1120
rect -4060 1058 -3579 1125
rect -4060 773 -3953 1058
rect -3657 773 -3579 1058
rect -4060 649 -3579 773
rect -4060 354 -3950 649
rect -3660 354 -3579 649
rect -3495 627 -3415 1177
rect -3272 1391 1400 1410
rect -3272 1236 -3225 1391
rect 1338 1236 1400 1391
rect -3272 959 1400 1236
rect -3272 627 -3196 959
rect -3495 420 -3196 627
rect 1313 492 1400 959
rect 1515 1193 2127 1410
rect 2347 1193 2697 1432
rect 1515 954 2697 1193
rect 1515 492 1610 954
rect 1313 420 1610 492
rect -3495 363 1610 420
rect -4060 197 -3579 354
rect -4427 -640 -4296 164
rect -4060 152 2291 197
rect 2374 188 2697 954
rect -4060 62 -3306 152
rect -4184 50 -3306 62
rect -4184 22 -3931 50
rect -4184 -246 -4107 22
rect -4183 -440 -4107 -246
rect -4427 -2024 -4406 -640
rect -4323 -2024 -4296 -640
rect -4186 -529 -4107 -440
rect -3997 -239 -3931 22
rect -3658 34 -3306 50
rect -3658 -239 -3513 34
rect -3997 -469 -3513 -239
rect -3399 -440 -3306 34
rect 1918 109 2291 152
rect 1918 -440 2440 109
rect -3399 -469 2440 -440
rect -3997 -518 2440 -469
rect -3997 -529 2439 -518
rect -4186 -555 2439 -529
rect -4186 -645 -3681 -555
rect 2244 -645 2439 -555
rect -4186 -680 2439 -645
rect -4427 -2590 -4296 -2024
rect -4427 -3616 -4395 -2590
rect -4321 -3616 -4296 -2590
rect -4175 -2108 -3937 -2103
rect -4175 -2142 2443 -2108
rect -4175 -2160 -3901 -2142
rect -4175 -3515 -4100 -2160
rect -4023 -2226 -3901 -2160
rect 2333 -2226 2443 -2142
rect -4023 -2259 2443 -2226
rect -4023 -3508 -3937 -2259
rect 2153 -2500 2443 -2259
rect 2153 -3508 2311 -2500
rect -4023 -3515 2311 -3508
rect -4175 -3535 2311 -3515
rect -4175 -3595 -3974 -3535
rect 2261 -3547 2311 -3535
rect 2378 -3547 2443 -2500
rect 2261 -3595 2443 -3547
rect -4175 -3606 2443 -3595
rect 2561 -2492 2697 188
rect 2561 -3189 2583 -2492
rect 2671 -3189 2697 -2492
rect 2561 -3231 2697 -3189
rect 2561 -3481 2574 -3231
rect 2685 -3481 2697 -3231
rect -4427 -3654 -4296 -3616
rect 2561 -3654 2697 -3481
rect -4427 -3672 2697 -3654
rect -4427 -3754 -4373 -3672
rect 2650 -3754 2697 -3672
rect -4427 -3755 2697 -3754
rect -4461 -3781 2731 -3755
rect -4461 -3815 -4401 -3781
rect 2671 -3815 2731 -3781
<< viali >>
rect -5024 -224 -4944 468
rect -4682 -92 -4602 600
rect -4332 6347 2644 6488
rect -4344 4172 -4257 6298
rect -4150 3889 2440 3929
rect -4064 1190 -3828 1431
rect -4349 1120 -4156 1182
rect -3415 627 -3272 1410
rect -3225 1236 1338 1391
rect 1400 492 1515 1410
rect 2127 1193 2347 1432
rect -4406 -2024 -4323 -640
rect -4107 -529 -3997 22
rect -3513 -469 -3399 34
rect -3681 -645 2244 -555
rect -4395 -3616 -4321 -2590
rect -4100 -3515 -4023 -2160
rect -3901 -2226 2333 -2142
rect -3974 -3595 2261 -3535
rect 2311 -3547 2378 -2500
rect 2583 -3189 2671 -2492
rect 2574 -3481 2685 -3231
rect -4373 -3754 2650 -3672
<< metal1 >>
rect -4365 6488 2686 6531
rect -4365 6347 -4332 6488
rect 2644 6347 2686 6488
rect -4365 6316 2686 6347
rect -4365 6298 -4234 6316
rect -4365 4172 -4344 6298
rect -4257 4172 -4234 6298
rect -4365 4140 -4234 4172
rect -4171 6114 2470 6178
rect -4171 5787 -4107 6114
rect -4072 5991 -4066 6055
rect -3950 5991 -3944 6055
rect -3756 5991 -3750 6055
rect -3634 5991 -3628 6055
rect -3440 5991 -3434 6055
rect -3318 5991 -3312 6055
rect -3124 5991 -3118 6055
rect -3002 5991 -2996 6055
rect -2808 5991 -2802 6055
rect -2686 5991 -2680 6055
rect -2492 5991 -2486 6055
rect -2370 5991 -2364 6055
rect -2176 5991 -2170 6055
rect -2054 5991 -2048 6055
rect -1860 5991 -1854 6055
rect -1738 5991 -1732 6055
rect -1544 5991 -1538 6055
rect -1422 5991 -1416 6055
rect -1228 5991 -1222 6055
rect -1106 5991 -1100 6055
rect -912 5991 -906 6055
rect -790 5991 -784 6055
rect -596 5991 -590 6055
rect -474 5991 -468 6055
rect -280 5991 -274 6055
rect -158 5991 -152 6055
rect 36 5991 42 6055
rect 158 5991 164 6055
rect 352 5991 358 6055
rect 474 5991 480 6055
rect 668 5991 674 6055
rect 790 5991 796 6055
rect 984 5991 990 6055
rect 1106 5991 1112 6055
rect 1300 5991 1306 6055
rect 1422 5991 1428 6055
rect 1616 5991 1622 6055
rect 1738 5991 1744 6055
rect 1932 5991 1938 6055
rect 2054 5991 2060 6055
rect 2248 5991 2254 6055
rect 2370 5991 2376 6055
rect -3914 5866 -3908 5930
rect -3792 5866 -3786 5930
rect -3598 5866 -3592 5930
rect -3476 5866 -3470 5930
rect -3282 5866 -3276 5930
rect -3160 5866 -3154 5930
rect -2966 5866 -2960 5930
rect -2844 5866 -2838 5930
rect -2650 5866 -2644 5930
rect -2528 5866 -2522 5930
rect -2334 5866 -2328 5930
rect -2212 5866 -2206 5930
rect -2018 5866 -2012 5930
rect -1896 5866 -1890 5930
rect -1702 5866 -1696 5930
rect -1580 5866 -1574 5930
rect -1386 5866 -1380 5930
rect -1264 5866 -1258 5930
rect -1070 5866 -1064 5930
rect -948 5866 -942 5930
rect -754 5866 -748 5930
rect -632 5866 -626 5930
rect -438 5866 -432 5930
rect -316 5866 -310 5930
rect -122 5866 -116 5930
rect 0 5866 6 5930
rect 194 5866 200 5930
rect 316 5866 322 5930
rect 510 5866 516 5930
rect 632 5866 638 5930
rect 826 5866 832 5930
rect 948 5866 954 5930
rect 1142 5866 1148 5930
rect 1264 5866 1270 5930
rect 1458 5866 1464 5930
rect 1580 5866 1586 5930
rect 1774 5866 1780 5930
rect 1896 5866 1902 5930
rect 2090 5866 2096 5930
rect 2212 5866 2218 5930
rect 2406 5787 2470 6114
rect -4171 5672 2470 5787
rect -4171 5360 -4107 5672
rect -4072 5551 -4066 5615
rect -3950 5551 -3944 5615
rect -3756 5551 -3750 5615
rect -3634 5551 -3628 5615
rect -3440 5551 -3434 5615
rect -3318 5551 -3312 5615
rect -3124 5551 -3118 5615
rect -3002 5551 -2996 5615
rect -2808 5551 -2802 5615
rect -2686 5551 -2680 5615
rect -2492 5551 -2486 5615
rect -2370 5551 -2364 5615
rect -2176 5551 -2170 5615
rect -2054 5551 -2048 5615
rect -1860 5551 -1854 5615
rect -1738 5551 -1732 5615
rect -1544 5551 -1538 5615
rect -1422 5551 -1416 5615
rect -1228 5551 -1222 5615
rect -1106 5551 -1100 5615
rect -912 5551 -906 5615
rect -790 5551 -784 5615
rect -596 5551 -590 5615
rect -474 5551 -468 5615
rect -280 5551 -274 5615
rect -158 5551 -152 5615
rect 36 5551 42 5615
rect 158 5551 164 5615
rect 352 5551 358 5615
rect 474 5551 480 5615
rect 668 5551 674 5615
rect 790 5551 796 5615
rect 984 5551 990 5615
rect 1106 5551 1112 5615
rect 1300 5551 1306 5615
rect 1422 5551 1428 5615
rect 1616 5551 1622 5615
rect 1738 5551 1744 5615
rect 1932 5551 1938 5615
rect 2054 5551 2060 5615
rect 2248 5551 2254 5615
rect 2370 5551 2376 5615
rect -3914 5426 -3908 5490
rect -3792 5426 -3786 5490
rect -3598 5426 -3592 5490
rect -3476 5426 -3470 5490
rect -3282 5426 -3276 5490
rect -3160 5426 -3154 5490
rect -2966 5426 -2960 5490
rect -2844 5426 -2838 5490
rect -2650 5426 -2644 5490
rect -2528 5426 -2522 5490
rect -2334 5426 -2328 5490
rect -2212 5426 -2206 5490
rect -2018 5426 -2012 5490
rect -1896 5426 -1890 5490
rect -1702 5426 -1696 5490
rect -1580 5426 -1574 5490
rect -1386 5426 -1380 5490
rect -1264 5426 -1258 5490
rect -1070 5426 -1064 5490
rect -948 5426 -942 5490
rect -754 5426 -748 5490
rect -632 5426 -626 5490
rect -438 5426 -432 5490
rect -316 5426 -310 5490
rect -122 5426 -116 5490
rect 0 5426 6 5490
rect 194 5426 200 5490
rect 316 5426 322 5490
rect 510 5426 516 5490
rect 632 5426 638 5490
rect 826 5426 832 5490
rect 948 5426 954 5490
rect 1142 5426 1148 5490
rect 1264 5426 1270 5490
rect 1458 5426 1464 5490
rect 1580 5426 1586 5490
rect 1774 5426 1780 5490
rect 1896 5426 1902 5490
rect 2090 5426 2096 5490
rect 2212 5426 2218 5490
rect 2406 5360 2470 5672
rect -4171 5245 2470 5360
rect -4171 4917 -4107 5245
rect -4072 5111 -4066 5175
rect -3950 5111 -3944 5175
rect -3756 5111 -3750 5175
rect -3634 5111 -3628 5175
rect -3440 5111 -3434 5175
rect -3318 5111 -3312 5175
rect -3124 5111 -3118 5175
rect -3002 5111 -2996 5175
rect -2808 5111 -2802 5175
rect -2686 5111 -2680 5175
rect -2492 5111 -2486 5175
rect -2370 5111 -2364 5175
rect -2176 5111 -2170 5175
rect -2054 5111 -2048 5175
rect -1860 5111 -1854 5175
rect -1738 5111 -1732 5175
rect -1544 5111 -1538 5175
rect -1422 5111 -1416 5175
rect -1228 5111 -1222 5175
rect -1106 5111 -1100 5175
rect -912 5111 -906 5175
rect -790 5111 -784 5175
rect -596 5111 -590 5175
rect -474 5111 -468 5175
rect -280 5111 -274 5175
rect -158 5111 -152 5175
rect 36 5111 42 5175
rect 158 5111 164 5175
rect 352 5111 358 5175
rect 474 5111 480 5175
rect 668 5111 674 5175
rect 790 5111 796 5175
rect 984 5111 990 5175
rect 1106 5111 1112 5175
rect 1300 5111 1306 5175
rect 1422 5111 1428 5175
rect 1616 5111 1622 5175
rect 1738 5111 1744 5175
rect 1932 5111 1938 5175
rect 2054 5111 2060 5175
rect 2248 5111 2254 5175
rect 2370 5111 2376 5175
rect -3914 4986 -3908 5050
rect -3792 4986 -3786 5050
rect -3598 4986 -3592 5050
rect -3476 4986 -3470 5050
rect -3282 4986 -3276 5050
rect -3160 4986 -3154 5050
rect -2966 4986 -2960 5050
rect -2844 4986 -2838 5050
rect -2650 4986 -2644 5050
rect -2528 4986 -2522 5050
rect -2334 4986 -2328 5050
rect -2212 4986 -2206 5050
rect -2018 4986 -2012 5050
rect -1896 4986 -1890 5050
rect -1702 4986 -1696 5050
rect -1580 4986 -1574 5050
rect -1386 4986 -1380 5050
rect -1264 4986 -1258 5050
rect -1070 4986 -1064 5050
rect -948 4986 -942 5050
rect -754 4986 -748 5050
rect -632 4986 -626 5050
rect -438 4986 -432 5050
rect -316 4986 -310 5050
rect -122 4986 -116 5050
rect 0 4986 6 5050
rect 194 4986 200 5050
rect 316 4986 322 5050
rect 510 4986 516 5050
rect 632 4986 638 5050
rect 826 4986 832 5050
rect 948 4986 954 5050
rect 1142 4986 1148 5050
rect 1264 4986 1270 5050
rect 1458 4986 1464 5050
rect 1580 4986 1586 5050
rect 1774 4986 1780 5050
rect 1896 4986 1902 5050
rect 2090 4986 2096 5050
rect 2212 4986 2218 5050
rect 2406 4917 2470 5245
rect -4171 4802 2470 4917
rect -4171 4484 -4107 4802
rect -4072 4676 -4066 4740
rect -3950 4676 -3944 4740
rect -3756 4676 -3750 4740
rect -3634 4676 -3628 4740
rect -3440 4676 -3434 4740
rect -3318 4676 -3312 4740
rect -3124 4676 -3118 4740
rect -3002 4676 -2996 4740
rect -2808 4676 -2802 4740
rect -2686 4676 -2680 4740
rect -2492 4676 -2486 4740
rect -2370 4676 -2364 4740
rect -2176 4676 -2170 4740
rect -2054 4676 -2048 4740
rect -1860 4676 -1854 4740
rect -1738 4676 -1732 4740
rect -1544 4676 -1538 4740
rect -1422 4676 -1416 4740
rect -1228 4676 -1222 4740
rect -1106 4676 -1100 4740
rect -912 4676 -906 4740
rect -790 4676 -784 4740
rect -596 4676 -590 4740
rect -474 4676 -468 4740
rect -280 4676 -274 4740
rect -158 4676 -152 4740
rect 36 4676 42 4740
rect 158 4676 164 4740
rect 352 4676 358 4740
rect 474 4676 480 4740
rect 668 4676 674 4740
rect 790 4676 796 4740
rect 984 4676 990 4740
rect 1106 4676 1112 4740
rect 1300 4676 1306 4740
rect 1422 4676 1428 4740
rect 1616 4676 1622 4740
rect 1738 4676 1744 4740
rect 1932 4676 1938 4740
rect 2054 4676 2060 4740
rect 2248 4676 2254 4740
rect 2370 4676 2376 4740
rect -3914 4551 -3908 4615
rect -3792 4551 -3786 4615
rect -3598 4551 -3592 4615
rect -3476 4551 -3470 4615
rect -3282 4551 -3276 4615
rect -3160 4551 -3154 4615
rect -2966 4551 -2960 4615
rect -2844 4551 -2838 4615
rect -2650 4551 -2644 4615
rect -2528 4551 -2522 4615
rect -2334 4551 -2328 4615
rect -2212 4551 -2206 4615
rect -2018 4551 -2012 4615
rect -1896 4551 -1890 4615
rect -1702 4551 -1696 4615
rect -1580 4551 -1574 4615
rect -1386 4551 -1380 4615
rect -1264 4551 -1258 4615
rect -1070 4551 -1064 4615
rect -948 4551 -942 4615
rect -754 4551 -748 4615
rect -632 4551 -626 4615
rect -438 4551 -432 4615
rect -316 4551 -310 4615
rect -122 4551 -116 4615
rect 0 4551 6 4615
rect 194 4551 200 4615
rect 316 4551 322 4615
rect 510 4551 516 4615
rect 632 4551 638 4615
rect 826 4551 832 4615
rect 948 4551 954 4615
rect 1142 4551 1148 4615
rect 1264 4551 1270 4615
rect 1458 4551 1464 4615
rect 1580 4551 1586 4615
rect 1774 4551 1780 4615
rect 1896 4551 1902 4615
rect 2090 4551 2096 4615
rect 2212 4551 2218 4615
rect 2406 4484 2470 4802
rect -4171 4369 2470 4484
rect -4171 4071 -4107 4369
rect -4072 4251 -4066 4315
rect -3950 4251 -3944 4315
rect -3756 4251 -3750 4315
rect -3634 4251 -3628 4315
rect -3440 4251 -3434 4315
rect -3318 4251 -3312 4315
rect -3124 4251 -3118 4315
rect -3002 4251 -2996 4315
rect -2808 4251 -2802 4315
rect -2686 4251 -2680 4315
rect -2492 4251 -2486 4315
rect -2370 4251 -2364 4315
rect -2176 4251 -2170 4315
rect -2054 4251 -2048 4315
rect -1860 4251 -1854 4315
rect -1738 4251 -1732 4315
rect -1544 4251 -1538 4315
rect -1422 4251 -1416 4315
rect -1228 4251 -1222 4315
rect -1106 4251 -1100 4315
rect -912 4251 -906 4315
rect -790 4251 -784 4315
rect -596 4251 -590 4315
rect -474 4251 -468 4315
rect -280 4251 -274 4315
rect -158 4251 -152 4315
rect 36 4251 42 4315
rect 158 4251 164 4315
rect 352 4251 358 4315
rect 474 4251 480 4315
rect 668 4251 674 4315
rect 790 4251 796 4315
rect 984 4251 990 4315
rect 1106 4251 1112 4315
rect 1300 4251 1306 4315
rect 1422 4251 1428 4315
rect 1616 4251 1622 4315
rect 1738 4251 1744 4315
rect 1932 4251 1938 4315
rect 2054 4251 2060 4315
rect 2248 4251 2254 4315
rect 2370 4251 2376 4315
rect -3914 4126 -3908 4190
rect -3792 4126 -3786 4190
rect -3598 4126 -3592 4190
rect -3476 4126 -3470 4190
rect -3282 4126 -3276 4190
rect -3160 4126 -3154 4190
rect -2966 4126 -2960 4190
rect -2844 4126 -2838 4190
rect -2650 4126 -2644 4190
rect -2528 4126 -2522 4190
rect -2334 4126 -2328 4190
rect -2212 4126 -2206 4190
rect -2018 4126 -2012 4190
rect -1896 4126 -1890 4190
rect -1702 4126 -1696 4190
rect -1580 4126 -1574 4190
rect -1386 4126 -1380 4190
rect -1264 4126 -1258 4190
rect -1070 4126 -1064 4190
rect -948 4126 -942 4190
rect -754 4126 -748 4190
rect -632 4126 -626 4190
rect -438 4126 -432 4190
rect -316 4126 -310 4190
rect -122 4126 -116 4190
rect 0 4126 6 4190
rect 194 4126 200 4190
rect 316 4126 322 4190
rect 510 4126 516 4190
rect 632 4126 638 4190
rect 826 4126 832 4190
rect 948 4126 954 4190
rect 1142 4126 1148 4190
rect 1264 4126 1270 4190
rect 1458 4126 1464 4190
rect 1580 4126 1586 4190
rect 1774 4126 1780 4190
rect 1896 4126 1902 4190
rect 2090 4126 2096 4190
rect 2212 4126 2218 4190
rect -4291 4066 -4107 4071
rect 2406 4066 2470 4369
rect -4291 4002 2470 4066
rect 2534 6106 2683 6131
rect -4291 1583 -4227 4002
rect -4170 3929 -4118 3941
rect 2350 3929 2485 3941
rect -4170 3889 -4150 3929
rect 2440 3889 2485 3929
rect -4170 3881 -4118 3889
rect 2350 3881 2485 3889
rect -4174 3757 2476 3821
rect -4174 3440 -4110 3757
rect -4072 3631 -4066 3695
rect -3950 3631 -3944 3695
rect -3756 3631 -3750 3695
rect -3634 3631 -3628 3695
rect -3440 3631 -3434 3695
rect -3318 3631 -3312 3695
rect -3124 3631 -3118 3695
rect -3002 3631 -2996 3695
rect -2808 3631 -2802 3695
rect -2686 3631 -2680 3695
rect -2492 3631 -2486 3695
rect -2370 3631 -2364 3695
rect -2176 3631 -2170 3695
rect -2054 3631 -2048 3695
rect -1860 3631 -1854 3695
rect -1738 3631 -1732 3695
rect -1544 3631 -1538 3695
rect -1422 3631 -1416 3695
rect -1228 3631 -1222 3695
rect -1106 3631 -1100 3695
rect -912 3631 -906 3695
rect -790 3631 -784 3695
rect -596 3631 -590 3695
rect -474 3631 -468 3695
rect -280 3631 -274 3695
rect -158 3631 -152 3695
rect 36 3631 42 3695
rect 158 3631 164 3695
rect 352 3631 358 3695
rect 474 3631 480 3695
rect 668 3631 674 3695
rect 790 3631 796 3695
rect 984 3631 990 3695
rect 1106 3631 1112 3695
rect 1300 3631 1306 3695
rect 1422 3631 1428 3695
rect 1616 3631 1622 3695
rect 1738 3631 1744 3695
rect 1932 3631 1938 3695
rect 2054 3631 2060 3695
rect 2248 3631 2254 3695
rect 2370 3631 2376 3695
rect -3914 3506 -3908 3570
rect -3792 3506 -3786 3570
rect -3598 3506 -3592 3570
rect -3476 3506 -3470 3570
rect -3282 3506 -3276 3570
rect -3160 3506 -3154 3570
rect -2966 3506 -2960 3570
rect -2844 3506 -2838 3570
rect -2650 3506 -2644 3570
rect -2528 3506 -2522 3570
rect -2334 3506 -2328 3570
rect -2212 3506 -2206 3570
rect -2018 3506 -2012 3570
rect -1896 3506 -1890 3570
rect -1702 3506 -1696 3570
rect -1580 3506 -1574 3570
rect -1386 3506 -1380 3570
rect -1264 3506 -1258 3570
rect -1070 3506 -1064 3570
rect -948 3506 -942 3570
rect -754 3506 -748 3570
rect -632 3506 -626 3570
rect -438 3506 -432 3570
rect -316 3506 -310 3570
rect -122 3506 -116 3570
rect 0 3506 6 3570
rect 194 3506 200 3570
rect 316 3506 322 3570
rect 510 3506 516 3570
rect 632 3506 638 3570
rect 826 3506 832 3570
rect 948 3506 954 3570
rect 1142 3506 1148 3570
rect 1264 3506 1270 3570
rect 1458 3506 1464 3570
rect 1580 3506 1586 3570
rect 1774 3506 1780 3570
rect 1896 3506 1902 3570
rect 2090 3506 2096 3570
rect 2212 3506 2218 3570
rect 2412 3440 2476 3757
rect -4174 3325 2476 3440
rect -4174 3002 -4110 3325
rect -4072 3196 -4066 3260
rect -3950 3196 -3944 3260
rect -3756 3196 -3750 3260
rect -3634 3196 -3628 3260
rect -3440 3196 -3434 3260
rect -3318 3196 -3312 3260
rect -3124 3196 -3118 3260
rect -3002 3196 -2996 3260
rect -2808 3196 -2802 3260
rect -2686 3196 -2680 3260
rect -2492 3196 -2486 3260
rect -2370 3196 -2364 3260
rect -2176 3196 -2170 3260
rect -2054 3196 -2048 3260
rect -1860 3196 -1854 3260
rect -1738 3196 -1732 3260
rect -1544 3196 -1538 3260
rect -1422 3196 -1416 3260
rect -1228 3196 -1222 3260
rect -1106 3196 -1100 3260
rect -912 3196 -906 3260
rect -790 3196 -784 3260
rect -596 3196 -590 3260
rect -474 3196 -468 3260
rect -280 3196 -274 3260
rect -158 3196 -152 3260
rect 36 3196 42 3260
rect 158 3196 164 3260
rect 352 3196 358 3260
rect 474 3196 480 3260
rect 668 3196 674 3260
rect 790 3196 796 3260
rect 984 3196 990 3260
rect 1106 3196 1112 3260
rect 1300 3196 1306 3260
rect 1422 3196 1428 3260
rect 1616 3196 1622 3260
rect 1738 3196 1744 3260
rect 1932 3196 1938 3260
rect 2054 3196 2060 3260
rect 2248 3196 2254 3260
rect 2370 3196 2376 3260
rect -3914 3071 -3908 3135
rect -3792 3071 -3786 3135
rect -3598 3071 -3592 3135
rect -3476 3071 -3470 3135
rect -3282 3071 -3276 3135
rect -3160 3071 -3154 3135
rect -2966 3071 -2960 3135
rect -2844 3071 -2838 3135
rect -2650 3071 -2644 3135
rect -2528 3071 -2522 3135
rect -2334 3071 -2328 3135
rect -2212 3071 -2206 3135
rect -2018 3071 -2012 3135
rect -1896 3071 -1890 3135
rect -1702 3071 -1696 3135
rect -1580 3071 -1574 3135
rect -1386 3071 -1380 3135
rect -1264 3071 -1258 3135
rect -1070 3071 -1064 3135
rect -948 3071 -942 3135
rect -754 3071 -748 3135
rect -632 3071 -626 3135
rect -438 3071 -432 3135
rect -316 3071 -310 3135
rect -122 3071 -116 3135
rect 0 3071 6 3135
rect 194 3071 200 3135
rect 316 3071 322 3135
rect 510 3071 516 3135
rect 632 3071 638 3135
rect 826 3071 832 3135
rect 948 3071 954 3135
rect 1142 3071 1148 3135
rect 1264 3071 1270 3135
rect 1458 3071 1464 3135
rect 1580 3071 1586 3135
rect 1774 3071 1780 3135
rect 1896 3071 1902 3135
rect 2090 3071 2096 3135
rect 2212 3071 2218 3135
rect 2412 3002 2476 3325
rect -4174 2887 2476 3002
rect -4174 2570 -4110 2887
rect -4072 2761 -4066 2825
rect -3950 2761 -3944 2825
rect -3756 2761 -3750 2825
rect -3634 2761 -3628 2825
rect -3440 2761 -3434 2825
rect -3318 2761 -3312 2825
rect -3124 2761 -3118 2825
rect -3002 2761 -2996 2825
rect -2808 2761 -2802 2825
rect -2686 2761 -2680 2825
rect -2492 2761 -2486 2825
rect -2370 2761 -2364 2825
rect -2176 2761 -2170 2825
rect -2054 2761 -2048 2825
rect -1860 2761 -1854 2825
rect -1738 2761 -1732 2825
rect -1544 2761 -1538 2825
rect -1422 2761 -1416 2825
rect -1228 2761 -1222 2825
rect -1106 2761 -1100 2825
rect -912 2761 -906 2825
rect -790 2761 -784 2825
rect -596 2761 -590 2825
rect -474 2761 -468 2825
rect -280 2761 -274 2825
rect -158 2761 -152 2825
rect 36 2761 42 2825
rect 158 2761 164 2825
rect 352 2761 358 2825
rect 474 2761 480 2825
rect 668 2761 674 2825
rect 790 2761 796 2825
rect 984 2761 990 2825
rect 1106 2761 1112 2825
rect 1300 2761 1306 2825
rect 1422 2761 1428 2825
rect 1616 2761 1622 2825
rect 1738 2761 1744 2825
rect 1932 2761 1938 2825
rect 2054 2761 2060 2825
rect 2248 2761 2254 2825
rect 2370 2761 2376 2825
rect -3914 2636 -3908 2700
rect -3792 2636 -3786 2700
rect -3598 2636 -3592 2700
rect -3476 2636 -3470 2700
rect -3282 2636 -3276 2700
rect -3160 2636 -3154 2700
rect -2966 2636 -2960 2700
rect -2844 2636 -2838 2700
rect -2650 2636 -2644 2700
rect -2528 2636 -2522 2700
rect -2334 2636 -2328 2700
rect -2212 2636 -2206 2700
rect -2018 2636 -2012 2700
rect -1896 2636 -1890 2700
rect -1702 2636 -1696 2700
rect -1580 2636 -1574 2700
rect -1386 2636 -1380 2700
rect -1264 2636 -1258 2700
rect -1070 2636 -1064 2700
rect -948 2636 -942 2700
rect -754 2636 -748 2700
rect -632 2636 -626 2700
rect -438 2636 -432 2700
rect -316 2636 -310 2700
rect -122 2636 -116 2700
rect 0 2636 6 2700
rect 194 2636 200 2700
rect 316 2636 322 2700
rect 510 2636 516 2700
rect 632 2636 638 2700
rect 826 2636 832 2700
rect 948 2636 954 2700
rect 1142 2636 1148 2700
rect 1264 2636 1270 2700
rect 1458 2636 1464 2700
rect 1580 2636 1586 2700
rect 1774 2636 1780 2700
rect 1896 2636 1902 2700
rect 2090 2636 2096 2700
rect 2212 2636 2218 2700
rect 2412 2570 2476 2887
rect -4174 2455 2476 2570
rect -4174 2135 -4110 2455
rect -4072 2326 -4066 2390
rect -3950 2326 -3944 2390
rect -3756 2326 -3750 2390
rect -3634 2326 -3628 2390
rect -3440 2326 -3434 2390
rect -3318 2326 -3312 2390
rect -3124 2326 -3118 2390
rect -3002 2326 -2996 2390
rect -2808 2326 -2802 2390
rect -2686 2326 -2680 2390
rect -2492 2326 -2486 2390
rect -2370 2326 -2364 2390
rect -2176 2326 -2170 2390
rect -2054 2326 -2048 2390
rect -1860 2326 -1854 2390
rect -1738 2326 -1732 2390
rect -1544 2326 -1538 2390
rect -1422 2326 -1416 2390
rect -1228 2326 -1222 2390
rect -1106 2326 -1100 2390
rect -912 2326 -906 2390
rect -790 2326 -784 2390
rect -596 2326 -590 2390
rect -474 2326 -468 2390
rect -280 2326 -274 2390
rect -158 2326 -152 2390
rect 36 2326 42 2390
rect 158 2326 164 2390
rect 352 2326 358 2390
rect 474 2326 480 2390
rect 668 2326 674 2390
rect 790 2326 796 2390
rect 984 2326 990 2390
rect 1106 2326 1112 2390
rect 1300 2326 1306 2390
rect 1422 2326 1428 2390
rect 1616 2326 1622 2390
rect 1738 2326 1744 2390
rect 1932 2326 1938 2390
rect 2054 2326 2060 2390
rect 2248 2326 2254 2390
rect 2370 2326 2376 2390
rect -3914 2201 -3908 2265
rect -3792 2201 -3786 2265
rect -3598 2201 -3592 2265
rect -3476 2201 -3470 2265
rect -3282 2201 -3276 2265
rect -3160 2201 -3154 2265
rect -2966 2201 -2960 2265
rect -2844 2201 -2838 2265
rect -2650 2201 -2644 2265
rect -2528 2201 -2522 2265
rect -2334 2201 -2328 2265
rect -2212 2201 -2206 2265
rect -2018 2201 -2012 2265
rect -1896 2201 -1890 2265
rect -1702 2201 -1696 2265
rect -1580 2201 -1574 2265
rect -1386 2201 -1380 2265
rect -1264 2201 -1258 2265
rect -1070 2201 -1064 2265
rect -948 2201 -942 2265
rect -754 2201 -748 2265
rect -632 2201 -626 2265
rect -438 2201 -432 2265
rect -316 2201 -310 2265
rect -122 2201 -116 2265
rect 0 2201 6 2265
rect 194 2201 200 2265
rect 316 2201 322 2265
rect 510 2201 516 2265
rect 632 2201 638 2265
rect 826 2201 832 2265
rect 948 2201 954 2265
rect 1142 2201 1148 2265
rect 1264 2201 1270 2265
rect 1458 2201 1464 2265
rect 1580 2201 1586 2265
rect 1774 2201 1780 2265
rect 1896 2201 1902 2265
rect 2090 2201 2096 2265
rect 2212 2201 2218 2265
rect 2412 2135 2476 2455
rect -4174 2040 2476 2135
rect -4174 1713 -4110 2040
rect -4072 1891 -4066 1955
rect -3950 1891 -3944 1955
rect -3756 1891 -3750 1955
rect -3634 1891 -3628 1955
rect -3440 1891 -3434 1955
rect -3318 1891 -3312 1955
rect -3124 1891 -3118 1955
rect -3002 1891 -2996 1955
rect -2808 1891 -2802 1955
rect -2686 1891 -2680 1955
rect -2492 1891 -2486 1955
rect -2370 1891 -2364 1955
rect -2176 1891 -2170 1955
rect -2054 1891 -2048 1955
rect -1860 1891 -1854 1955
rect -1738 1891 -1732 1955
rect -1544 1891 -1538 1955
rect -1422 1891 -1416 1955
rect -1228 1891 -1222 1955
rect -1106 1891 -1100 1955
rect -912 1891 -906 1955
rect -790 1891 -784 1955
rect -596 1891 -590 1955
rect -474 1891 -468 1955
rect -280 1891 -274 1955
rect -158 1891 -152 1955
rect 36 1891 42 1955
rect 158 1891 164 1955
rect 352 1891 358 1955
rect 474 1891 480 1955
rect 668 1891 674 1955
rect 790 1891 796 1955
rect 984 1891 990 1955
rect 1106 1891 1112 1955
rect 1300 1891 1306 1955
rect 1422 1891 1428 1955
rect 1616 1891 1622 1955
rect 1738 1891 1744 1955
rect 1932 1891 1938 1955
rect 2054 1891 2060 1955
rect 2248 1891 2254 1955
rect 2370 1891 2376 1955
rect -3914 1766 -3908 1830
rect -3792 1766 -3786 1830
rect -3598 1766 -3592 1830
rect -3476 1766 -3470 1830
rect -3282 1766 -3276 1830
rect -3160 1766 -3154 1830
rect -2966 1766 -2960 1830
rect -2844 1766 -2838 1830
rect -2650 1766 -2644 1830
rect -2528 1766 -2522 1830
rect -2334 1766 -2328 1830
rect -2212 1766 -2206 1830
rect -2018 1766 -2012 1830
rect -1896 1766 -1890 1830
rect -1702 1766 -1696 1830
rect -1580 1766 -1574 1830
rect -1386 1766 -1380 1830
rect -1264 1766 -1258 1830
rect -1070 1766 -1064 1830
rect -948 1766 -942 1830
rect -754 1766 -748 1830
rect -632 1766 -626 1830
rect -438 1766 -432 1830
rect -316 1766 -310 1830
rect -122 1766 -116 1830
rect 0 1766 6 1830
rect 194 1766 200 1830
rect 316 1766 322 1830
rect 510 1766 516 1830
rect 632 1766 638 1830
rect 826 1766 832 1830
rect 948 1766 954 1830
rect 1142 1766 1148 1830
rect 1264 1766 1270 1830
rect 1458 1766 1464 1830
rect 1580 1766 1586 1830
rect 1774 1766 1780 1830
rect 1896 1766 1902 1830
rect 2090 1766 2096 1830
rect 2212 1766 2218 1830
rect 2412 1713 2476 2040
rect -4174 1649 2476 1713
rect -4291 1519 -3634 1583
rect 2412 1569 2476 1649
rect -4077 1431 -3813 1445
rect -4362 1182 -4140 1401
rect -4362 1120 -4349 1182
rect -4156 1120 -4140 1182
rect -4077 1190 -4064 1431
rect -3828 1190 -3813 1431
rect -4077 1177 -3813 1190
rect -4362 1106 -4140 1120
rect -4361 950 -4126 1019
rect -4862 858 -4126 950
rect -4858 722 -4744 858
rect -4361 819 -4126 858
rect -3826 819 -3808 1019
rect -5004 480 -4994 578
rect -5030 468 -4994 480
rect -5030 -224 -5024 468
rect -4930 -14 -4920 578
rect -4838 340 -4766 722
rect -4688 600 -4596 612
rect -4688 572 -4682 600
rect -4944 -224 -4938 -14
rect -4844 -194 -4772 170
rect -4690 -10 -4682 572
rect -4688 -92 -4682 -10
rect -4602 -92 -4596 600
rect -4361 489 -4126 689
rect -3826 489 -3762 689
rect -3846 452 -3762 489
rect -3698 491 -3634 1519
rect 1911 1506 2476 1569
rect 1911 1505 2412 1506
rect -3444 1426 1553 1449
rect -3444 1410 -3185 1426
rect -3444 627 -3415 1410
rect -3272 1391 -3185 1410
rect 1307 1410 1553 1426
rect 1307 1391 1400 1410
rect -3272 1236 -3225 1391
rect 1338 1236 1400 1391
rect -3272 1196 -3185 1236
rect 1307 1196 1400 1236
rect -3272 1181 1400 1196
rect -3272 627 -3246 1181
rect -2947 1177 -1099 1181
rect 447 1177 749 1181
rect -3444 598 -3246 627
rect -3113 596 -3064 840
rect -2947 640 -2854 1177
rect -2746 874 -2386 911
rect -2746 596 -2697 874
rect -3113 560 -2697 596
rect -3113 506 -3064 560
rect -2746 506 -2697 560
rect -2529 507 -2480 840
rect -2423 595 -2386 874
rect -2356 638 -2263 1177
rect -2424 559 -2217 595
rect -2159 507 -2110 840
rect -3698 436 -3438 491
rect -3269 436 -3262 491
rect -3113 424 -2697 506
rect -2595 491 -2110 507
rect -2595 436 -2531 491
rect -3113 423 -2701 424
rect -4361 325 -4126 364
rect -4361 244 -3762 325
rect -4361 164 -4126 244
rect -3846 167 -3762 244
rect -3228 227 -3222 279
rect -3081 227 -3075 279
rect -4688 -104 -4596 -92
rect -4392 22 -3980 34
rect -4392 2 -4107 22
rect -5030 -236 -4938 -224
rect -4864 -348 -4750 -194
rect -4392 -308 -4373 2
rect -4134 -308 -4107 2
rect -4892 -438 -4882 -348
rect -4728 -372 -4718 -348
rect -4392 -372 -4107 -308
rect -4728 -438 -4107 -372
rect -4862 -458 -4107 -438
rect -4392 -529 -4107 -458
rect -3997 -198 -3980 22
rect -3846 22 -3829 167
rect -3774 22 -3762 167
rect -3846 -143 -3762 22
rect -3537 34 -3380 56
rect -3537 -198 -3513 34
rect -3997 -335 -3513 -198
rect -3997 -529 -3980 -335
rect -3909 -469 -3892 -408
rect -3713 -469 -3702 -408
rect -3537 -469 -3513 -335
rect -3399 -469 -3380 34
rect -3221 -69 -3156 -60
rect -3221 -250 -3214 -69
rect -3162 -250 -3156 -69
rect -3221 -256 -3156 -250
rect -3123 -329 -3084 227
rect -3028 -253 -2937 423
rect -2595 421 -2110 436
rect -1946 595 -1897 840
rect -1779 636 -1686 1177
rect -1578 878 -1220 915
rect -1578 595 -1529 878
rect -1946 559 -1529 595
rect -1946 504 -1897 559
rect -1578 504 -1529 559
rect -1946 423 -1529 504
rect -1356 504 -1307 840
rect -1257 595 -1220 878
rect -1192 638 -1099 1177
rect -1263 559 -1056 595
rect -996 504 -947 840
rect -1356 489 -947 504
rect -2795 323 -2789 375
rect -2648 323 -2642 375
rect -2788 -69 -2723 -60
rect -2788 -250 -2776 -69
rect -2724 -250 -2723 -69
rect -2788 -256 -2723 -250
rect -2693 -322 -2653 323
rect -2595 -256 -2505 421
rect -1927 227 -1921 279
rect -1780 227 -1774 279
rect -2284 80 -2192 86
rect -2284 20 -2192 28
rect -4392 -546 -3980 -529
rect -4392 -547 -4120 -546
rect -4434 -640 -4296 -607
rect -3892 -621 -3825 -469
rect -3537 -486 -3380 -469
rect -2407 -531 -2312 -58
rect -2256 -316 -2214 20
rect -2183 -66 -2118 -60
rect -2183 -247 -2178 -66
rect -2126 -247 -2118 -66
rect -2183 -256 -2118 -247
rect -1916 -67 -1851 -60
rect -1916 -248 -1907 -67
rect -1855 -248 -1851 -67
rect -1916 -256 -1851 -248
rect -1822 -329 -1781 227
rect -1724 -253 -1639 423
rect -1356 422 -947 434
rect -1495 323 -1489 375
rect -1348 323 -1342 375
rect -1485 -66 -1420 -60
rect -1485 -247 -1478 -66
rect -1426 -247 -1420 -66
rect -1485 -256 -1420 -247
rect -1389 -320 -1350 323
rect -1290 -256 -1199 422
rect -779 153 -733 840
rect -622 836 -510 848
rect -622 648 -611 836
rect -520 648 -510 836
rect -622 638 -510 648
rect -665 375 -624 585
rect -502 375 -461 581
rect -665 323 -657 375
rect -470 323 -461 375
rect -410 153 -364 840
rect -981 80 -889 86
rect -779 54 -364 153
rect -191 152 -145 840
rect -36 834 76 847
rect -36 646 -26 834
rect 65 646 76 834
rect -36 637 76 646
rect -85 279 -44 580
rect 74 279 115 582
rect -86 227 -79 279
rect 108 227 116 279
rect 185 152 231 840
rect 388 834 500 846
rect 388 646 396 834
rect 487 646 500 834
rect 388 636 500 646
rect 539 640 667 1177
rect 707 837 819 849
rect 707 649 716 837
rect 807 649 819 837
rect 986 822 1073 828
rect 1072 659 1073 822
rect 986 652 1073 659
rect 707 639 819 649
rect 1168 599 1202 844
rect 1059 598 1202 599
rect 479 555 1202 598
rect 1059 551 1202 555
rect -981 20 -889 28
rect -1108 -531 -1013 -54
rect -955 -318 -913 20
rect -881 -66 -816 -60
rect -881 -247 -874 -66
rect -822 -247 -816 -66
rect -881 -256 -816 -247
rect -685 -408 -580 54
rect -191 51 231 152
rect 10 13 122 51
rect -475 6 122 13
rect -523 -21 122 6
rect 325 -19 1114 16
rect -523 -317 -484 -21
rect -402 -255 -136 -59
rect -720 -469 -713 -408
rect -559 -469 -551 -408
rect -341 -531 -206 -255
rect -87 -317 -48 -21
rect 10 -257 122 -21
rect 402 -65 484 -57
rect 244 -85 326 -78
rect 244 -254 250 -85
rect 317 -254 326 -85
rect 402 -234 408 -65
rect 475 -234 484 -65
rect 719 -65 801 -56
rect 402 -241 484 -234
rect 563 -83 645 -76
rect 244 -262 326 -254
rect 563 -252 569 -83
rect 636 -252 645 -83
rect 719 -234 725 -65
rect 792 -234 801 -65
rect 719 -240 801 -234
rect 879 -82 961 -74
rect 563 -260 645 -252
rect 879 -251 887 -82
rect 954 -251 961 -82
rect 879 -258 961 -251
rect 1028 -78 1114 -19
rect 1028 -255 1035 -78
rect 1107 -255 1114 -78
rect 1028 -302 1114 -255
rect 1159 -257 1197 551
rect 1373 492 1400 1181
rect 1515 492 1553 1410
rect 1373 461 1553 492
rect 1911 489 1975 1505
rect 2534 1495 2683 1506
rect 1716 434 1725 489
rect 1966 434 1975 489
rect 2111 1432 2683 1445
rect 2111 1193 2127 1432
rect 2347 1193 2683 1432
rect 2111 1091 2683 1193
rect 1693 174 1726 175
rect 1583 122 1589 174
rect 1726 122 1732 174
rect 1458 70 1529 78
rect 1231 -15 1458 15
rect 1312 -80 1394 -72
rect 1312 -249 1320 -80
rect 1387 -249 1394 -80
rect 1312 -256 1394 -249
rect 320 -324 1458 -302
rect 1529 -186 1616 -123
rect 1693 -308 1726 122
rect 320 -332 1529 -324
rect 1790 -367 1841 -54
rect 2111 -213 2363 1091
rect 2453 1015 2683 1026
rect 2453 681 2534 1015
rect 2453 616 2683 681
rect 2453 126 2683 381
rect 2453 -122 2683 -109
rect 2111 -283 2699 -213
rect 1790 -437 2589 -367
rect -4434 -2024 -4406 -640
rect -4323 -2024 -4296 -640
rect -4196 -688 -3825 -621
rect -3707 -555 2271 -531
rect -3707 -645 -3681 -555
rect 2244 -645 2271 -555
rect -3707 -660 2271 -645
rect -4196 -756 -4129 -688
rect -4196 -823 2475 -756
rect -4196 -1125 -4129 -823
rect -4072 -942 -4066 -878
rect -3950 -942 -3944 -878
rect -3756 -942 -3750 -878
rect -3634 -942 -3628 -878
rect -3440 -942 -3434 -878
rect -3318 -942 -3312 -878
rect -3124 -942 -3118 -878
rect -3002 -942 -2996 -878
rect -2808 -942 -2802 -878
rect -2686 -942 -2680 -878
rect -2492 -942 -2486 -878
rect -2370 -942 -2364 -878
rect -2176 -942 -2170 -878
rect -2054 -942 -2048 -878
rect -1860 -942 -1854 -878
rect -1738 -942 -1732 -878
rect -1544 -942 -1538 -878
rect -1422 -942 -1416 -878
rect -1228 -942 -1222 -878
rect -1106 -942 -1100 -878
rect -912 -942 -906 -878
rect -790 -942 -784 -878
rect -596 -942 -590 -878
rect -474 -942 -468 -878
rect -280 -942 -274 -878
rect -158 -942 -152 -878
rect 36 -942 42 -878
rect 158 -942 164 -878
rect 352 -942 358 -878
rect 474 -942 480 -878
rect 668 -942 674 -878
rect 790 -942 796 -878
rect 984 -942 990 -878
rect 1106 -942 1112 -878
rect 1300 -942 1306 -878
rect 1422 -942 1428 -878
rect 1616 -942 1622 -878
rect 1738 -942 1744 -878
rect 1932 -942 1938 -878
rect 2054 -942 2060 -878
rect 2248 -942 2254 -878
rect 2370 -942 2376 -878
rect -3914 -1067 -3908 -1003
rect -3792 -1067 -3786 -1003
rect -3598 -1067 -3592 -1003
rect -3476 -1067 -3470 -1003
rect -3282 -1067 -3276 -1003
rect -3160 -1067 -3154 -1003
rect -2966 -1067 -2960 -1003
rect -2844 -1067 -2838 -1003
rect -2650 -1067 -2644 -1003
rect -2528 -1067 -2522 -1003
rect -2334 -1067 -2328 -1003
rect -2212 -1067 -2206 -1003
rect -2018 -1067 -2012 -1003
rect -1896 -1067 -1890 -1003
rect -1702 -1067 -1696 -1003
rect -1580 -1067 -1574 -1003
rect -1386 -1067 -1380 -1003
rect -1264 -1067 -1258 -1003
rect -1070 -1067 -1064 -1003
rect -948 -1067 -942 -1003
rect -754 -1067 -748 -1003
rect -632 -1067 -626 -1003
rect -438 -1067 -432 -1003
rect -316 -1067 -310 -1003
rect -122 -1067 -116 -1003
rect 0 -1067 6 -1003
rect 194 -1067 200 -1003
rect 316 -1067 322 -1003
rect 510 -1067 516 -1003
rect 632 -1067 638 -1003
rect 826 -1067 832 -1003
rect 948 -1067 954 -1003
rect 1142 -1067 1148 -1003
rect 1264 -1067 1270 -1003
rect 1458 -1067 1464 -1003
rect 1580 -1067 1586 -1003
rect 1774 -1067 1780 -1003
rect 1896 -1067 1902 -1003
rect 2090 -1067 2096 -1003
rect 2212 -1067 2218 -1003
rect 2408 -1125 2475 -823
rect -4196 -1240 2475 -1125
rect -4196 -1546 -4129 -1240
rect -4072 -1360 -4066 -1296
rect -3950 -1360 -3944 -1296
rect -3756 -1360 -3750 -1296
rect -3634 -1360 -3628 -1296
rect -3440 -1360 -3434 -1296
rect -3318 -1360 -3312 -1296
rect -3124 -1360 -3118 -1296
rect -3002 -1360 -2996 -1296
rect -2808 -1360 -2802 -1296
rect -2686 -1360 -2680 -1296
rect -2492 -1360 -2486 -1296
rect -2370 -1360 -2364 -1296
rect -2176 -1360 -2170 -1296
rect -2054 -1360 -2048 -1296
rect -1860 -1360 -1854 -1296
rect -1738 -1360 -1732 -1296
rect -1544 -1360 -1538 -1296
rect -1422 -1360 -1416 -1296
rect -1228 -1360 -1222 -1296
rect -1106 -1360 -1100 -1296
rect -912 -1360 -906 -1296
rect -790 -1360 -784 -1296
rect -596 -1360 -590 -1296
rect -474 -1360 -468 -1296
rect -280 -1360 -274 -1296
rect -158 -1360 -152 -1296
rect 36 -1360 42 -1296
rect 158 -1360 164 -1296
rect 352 -1360 358 -1296
rect 474 -1360 480 -1296
rect 668 -1360 674 -1296
rect 790 -1360 796 -1296
rect 984 -1360 990 -1296
rect 1106 -1360 1112 -1296
rect 1300 -1360 1306 -1296
rect 1422 -1360 1428 -1296
rect 1616 -1360 1622 -1296
rect 1738 -1360 1744 -1296
rect 1932 -1360 1938 -1296
rect 2054 -1360 2060 -1296
rect 2248 -1360 2254 -1296
rect 2370 -1360 2376 -1296
rect -3914 -1485 -3908 -1421
rect -3792 -1485 -3786 -1421
rect -3598 -1485 -3592 -1421
rect -3476 -1485 -3470 -1421
rect -3282 -1485 -3276 -1421
rect -3160 -1485 -3154 -1421
rect -2966 -1485 -2960 -1421
rect -2844 -1485 -2838 -1421
rect -2650 -1485 -2644 -1421
rect -2528 -1485 -2522 -1421
rect -2334 -1485 -2328 -1421
rect -2212 -1485 -2206 -1421
rect -2018 -1485 -2012 -1421
rect -1896 -1485 -1890 -1421
rect -1702 -1485 -1696 -1421
rect -1580 -1485 -1574 -1421
rect -1386 -1485 -1380 -1421
rect -1264 -1485 -1258 -1421
rect -1070 -1485 -1064 -1421
rect -948 -1485 -942 -1421
rect -754 -1485 -748 -1421
rect -632 -1485 -626 -1421
rect -438 -1485 -432 -1421
rect -316 -1485 -310 -1421
rect -122 -1485 -116 -1421
rect 0 -1485 6 -1421
rect 194 -1485 200 -1421
rect 316 -1485 322 -1421
rect 510 -1485 516 -1421
rect 632 -1485 638 -1421
rect 826 -1485 832 -1421
rect 948 -1485 954 -1421
rect 1142 -1485 1148 -1421
rect 1264 -1485 1270 -1421
rect 1458 -1485 1464 -1421
rect 1580 -1485 1586 -1421
rect 1774 -1485 1780 -1421
rect 1896 -1485 1902 -1421
rect 2090 -1485 2096 -1421
rect 2212 -1485 2218 -1421
rect 2408 -1546 2475 -1240
rect -4196 -1661 2475 -1546
rect -4196 -1956 -4129 -1661
rect -4072 -1778 -4066 -1714
rect -3950 -1778 -3944 -1714
rect -3756 -1778 -3750 -1714
rect -3634 -1778 -3628 -1714
rect -3440 -1778 -3434 -1714
rect -3318 -1778 -3312 -1714
rect -3124 -1778 -3118 -1714
rect -3002 -1778 -2996 -1714
rect -2808 -1778 -2802 -1714
rect -2686 -1778 -2680 -1714
rect -2492 -1778 -2486 -1714
rect -2370 -1778 -2364 -1714
rect -2176 -1778 -2170 -1714
rect -2054 -1778 -2048 -1714
rect -1860 -1778 -1854 -1714
rect -1738 -1778 -1732 -1714
rect -1544 -1778 -1538 -1714
rect -1422 -1778 -1416 -1714
rect -1228 -1778 -1222 -1714
rect -1106 -1778 -1100 -1714
rect -912 -1778 -906 -1714
rect -790 -1778 -784 -1714
rect -596 -1778 -590 -1714
rect -474 -1778 -468 -1714
rect -280 -1778 -274 -1714
rect -158 -1778 -152 -1714
rect 36 -1778 42 -1714
rect 158 -1778 164 -1714
rect 352 -1778 358 -1714
rect 474 -1778 480 -1714
rect 668 -1778 674 -1714
rect 790 -1778 796 -1714
rect 984 -1778 990 -1714
rect 1106 -1778 1112 -1714
rect 1300 -1778 1306 -1714
rect 1422 -1778 1428 -1714
rect 1616 -1778 1622 -1714
rect 1738 -1778 1744 -1714
rect 1932 -1778 1938 -1714
rect 2054 -1778 2060 -1714
rect 2248 -1778 2254 -1714
rect 2370 -1778 2376 -1714
rect -3914 -1903 -3908 -1839
rect -3792 -1903 -3786 -1839
rect -3598 -1903 -3592 -1839
rect -3476 -1903 -3470 -1839
rect -3282 -1903 -3276 -1839
rect -3160 -1903 -3154 -1839
rect -2966 -1903 -2960 -1839
rect -2844 -1903 -2838 -1839
rect -2650 -1903 -2644 -1839
rect -2528 -1903 -2522 -1839
rect -2334 -1903 -2328 -1839
rect -2212 -1903 -2206 -1839
rect -2018 -1903 -2012 -1839
rect -1896 -1903 -1890 -1839
rect -1702 -1903 -1696 -1839
rect -1580 -1903 -1574 -1839
rect -1386 -1903 -1380 -1839
rect -1264 -1903 -1258 -1839
rect -1070 -1903 -1064 -1839
rect -948 -1903 -942 -1839
rect -754 -1903 -748 -1839
rect -632 -1903 -626 -1839
rect -438 -1903 -432 -1839
rect -316 -1903 -310 -1839
rect -122 -1903 -116 -1839
rect 0 -1903 6 -1839
rect 194 -1903 200 -1839
rect 316 -1903 322 -1839
rect 510 -1903 516 -1839
rect 632 -1903 638 -1839
rect 826 -1903 832 -1839
rect 948 -1903 954 -1839
rect 1142 -1903 1148 -1839
rect 1264 -1903 1270 -1839
rect 1458 -1903 1464 -1839
rect 1580 -1903 1586 -1839
rect 1774 -1903 1780 -1839
rect 1896 -1903 1902 -1839
rect 2090 -1903 2096 -1839
rect 2212 -1903 2218 -1839
rect 2408 -1956 2475 -1661
rect -4196 -2023 2475 -1956
rect -4434 -2055 -4296 -2024
rect -4392 -2110 2353 -2099
rect -4392 -2460 -4382 -2110
rect -4133 -2142 2353 -2110
rect -4133 -2160 -3901 -2142
rect -4133 -2460 -4100 -2160
rect -4392 -2472 -4100 -2460
rect -4434 -2590 -4296 -2548
rect -4434 -3616 -4395 -2590
rect -4321 -3616 -4296 -2590
rect -4125 -3515 -4100 -2472
rect -4023 -2226 -3901 -2160
rect 2333 -2226 2353 -2142
rect -4023 -2255 2353 -2226
rect -4023 -3515 -3994 -2255
rect -3792 -2735 -3434 -2402
rect -3792 -3361 -3434 -3028
rect -3253 -3372 -3053 -2255
rect -4125 -3517 -3994 -3515
rect -2853 -3517 -2653 -2426
rect -2453 -3372 -2253 -2255
rect -2053 -3517 -1853 -2426
rect -1653 -3372 -1453 -2255
rect -1253 -3517 -1053 -2426
rect -853 -3372 -653 -2255
rect -453 -3517 -253 -2426
rect -53 -3372 147 -2255
rect 347 -3517 547 -2426
rect 747 -3372 947 -2255
rect 2519 -2364 2589 -437
rect 1147 -3517 1347 -2426
rect 1604 -2434 2589 -2364
rect 2629 -2469 2699 -283
rect 2290 -2500 2402 -2478
rect 1621 -3043 1979 -2710
rect 1598 -3267 2228 -3239
rect 1598 -3441 1627 -3267
rect 2200 -3441 2228 -3267
rect 1598 -3466 2228 -3441
rect 2290 -3517 2311 -2500
rect -4125 -3535 2311 -3517
rect -4125 -3595 -3974 -3535
rect 2261 -3547 2311 -3535
rect 2378 -3547 2402 -2500
rect 2261 -3595 2402 -3547
rect -4125 -3606 2402 -3595
rect 2561 -2492 2699 -2469
rect 2561 -3189 2583 -2492
rect 2671 -3189 2699 -2492
rect 2561 -3220 2699 -3189
rect 2561 -3231 2629 -3220
rect 2561 -3481 2574 -3231
rect 2561 -3491 2629 -3481
rect -4434 -3654 -4296 -3616
rect 2561 -3654 2699 -3491
rect -4434 -3672 2699 -3654
rect -4434 -3754 -4373 -3672
rect 2650 -3754 2699 -3672
rect -4434 -3792 2699 -3754
<< via1 >>
rect -4332 6347 2644 6488
rect -4066 5991 -3950 6055
rect -3750 5991 -3634 6055
rect -3434 5991 -3318 6055
rect -3118 5991 -3002 6055
rect -2802 5991 -2686 6055
rect -2486 5991 -2370 6055
rect -2170 5991 -2054 6055
rect -1854 5991 -1738 6055
rect -1538 5991 -1422 6055
rect -1222 5991 -1106 6055
rect -906 5991 -790 6055
rect -590 5991 -474 6055
rect -274 5991 -158 6055
rect 42 5991 158 6055
rect 358 5991 474 6055
rect 674 5991 790 6055
rect 990 5991 1106 6055
rect 1306 5991 1422 6055
rect 1622 5991 1738 6055
rect 1938 5991 2054 6055
rect 2254 5991 2370 6055
rect -3908 5866 -3792 5930
rect -3592 5866 -3476 5930
rect -3276 5866 -3160 5930
rect -2960 5866 -2844 5930
rect -2644 5866 -2528 5930
rect -2328 5866 -2212 5930
rect -2012 5866 -1896 5930
rect -1696 5866 -1580 5930
rect -1380 5866 -1264 5930
rect -1064 5866 -948 5930
rect -748 5866 -632 5930
rect -432 5866 -316 5930
rect -116 5866 0 5930
rect 200 5866 316 5930
rect 516 5866 632 5930
rect 832 5866 948 5930
rect 1148 5866 1264 5930
rect 1464 5866 1580 5930
rect 1780 5866 1896 5930
rect 2096 5866 2212 5930
rect -4066 5551 -3950 5615
rect -3750 5551 -3634 5615
rect -3434 5551 -3318 5615
rect -3118 5551 -3002 5615
rect -2802 5551 -2686 5615
rect -2486 5551 -2370 5615
rect -2170 5551 -2054 5615
rect -1854 5551 -1738 5615
rect -1538 5551 -1422 5615
rect -1222 5551 -1106 5615
rect -906 5551 -790 5615
rect -590 5551 -474 5615
rect -274 5551 -158 5615
rect 42 5551 158 5615
rect 358 5551 474 5615
rect 674 5551 790 5615
rect 990 5551 1106 5615
rect 1306 5551 1422 5615
rect 1622 5551 1738 5615
rect 1938 5551 2054 5615
rect 2254 5551 2370 5615
rect -3908 5426 -3792 5490
rect -3592 5426 -3476 5490
rect -3276 5426 -3160 5490
rect -2960 5426 -2844 5490
rect -2644 5426 -2528 5490
rect -2328 5426 -2212 5490
rect -2012 5426 -1896 5490
rect -1696 5426 -1580 5490
rect -1380 5426 -1264 5490
rect -1064 5426 -948 5490
rect -748 5426 -632 5490
rect -432 5426 -316 5490
rect -116 5426 0 5490
rect 200 5426 316 5490
rect 516 5426 632 5490
rect 832 5426 948 5490
rect 1148 5426 1264 5490
rect 1464 5426 1580 5490
rect 1780 5426 1896 5490
rect 2096 5426 2212 5490
rect -4066 5111 -3950 5175
rect -3750 5111 -3634 5175
rect -3434 5111 -3318 5175
rect -3118 5111 -3002 5175
rect -2802 5111 -2686 5175
rect -2486 5111 -2370 5175
rect -2170 5111 -2054 5175
rect -1854 5111 -1738 5175
rect -1538 5111 -1422 5175
rect -1222 5111 -1106 5175
rect -906 5111 -790 5175
rect -590 5111 -474 5175
rect -274 5111 -158 5175
rect 42 5111 158 5175
rect 358 5111 474 5175
rect 674 5111 790 5175
rect 990 5111 1106 5175
rect 1306 5111 1422 5175
rect 1622 5111 1738 5175
rect 1938 5111 2054 5175
rect 2254 5111 2370 5175
rect -3908 4986 -3792 5050
rect -3592 4986 -3476 5050
rect -3276 4986 -3160 5050
rect -2960 4986 -2844 5050
rect -2644 4986 -2528 5050
rect -2328 4986 -2212 5050
rect -2012 4986 -1896 5050
rect -1696 4986 -1580 5050
rect -1380 4986 -1264 5050
rect -1064 4986 -948 5050
rect -748 4986 -632 5050
rect -432 4986 -316 5050
rect -116 4986 0 5050
rect 200 4986 316 5050
rect 516 4986 632 5050
rect 832 4986 948 5050
rect 1148 4986 1264 5050
rect 1464 4986 1580 5050
rect 1780 4986 1896 5050
rect 2096 4986 2212 5050
rect -4066 4676 -3950 4740
rect -3750 4676 -3634 4740
rect -3434 4676 -3318 4740
rect -3118 4676 -3002 4740
rect -2802 4676 -2686 4740
rect -2486 4676 -2370 4740
rect -2170 4676 -2054 4740
rect -1854 4676 -1738 4740
rect -1538 4676 -1422 4740
rect -1222 4676 -1106 4740
rect -906 4676 -790 4740
rect -590 4676 -474 4740
rect -274 4676 -158 4740
rect 42 4676 158 4740
rect 358 4676 474 4740
rect 674 4676 790 4740
rect 990 4676 1106 4740
rect 1306 4676 1422 4740
rect 1622 4676 1738 4740
rect 1938 4676 2054 4740
rect 2254 4676 2370 4740
rect -3908 4551 -3792 4615
rect -3592 4551 -3476 4615
rect -3276 4551 -3160 4615
rect -2960 4551 -2844 4615
rect -2644 4551 -2528 4615
rect -2328 4551 -2212 4615
rect -2012 4551 -1896 4615
rect -1696 4551 -1580 4615
rect -1380 4551 -1264 4615
rect -1064 4551 -948 4615
rect -748 4551 -632 4615
rect -432 4551 -316 4615
rect -116 4551 0 4615
rect 200 4551 316 4615
rect 516 4551 632 4615
rect 832 4551 948 4615
rect 1148 4551 1264 4615
rect 1464 4551 1580 4615
rect 1780 4551 1896 4615
rect 2096 4551 2212 4615
rect -4066 4251 -3950 4315
rect -3750 4251 -3634 4315
rect -3434 4251 -3318 4315
rect -3118 4251 -3002 4315
rect -2802 4251 -2686 4315
rect -2486 4251 -2370 4315
rect -2170 4251 -2054 4315
rect -1854 4251 -1738 4315
rect -1538 4251 -1422 4315
rect -1222 4251 -1106 4315
rect -906 4251 -790 4315
rect -590 4251 -474 4315
rect -274 4251 -158 4315
rect 42 4251 158 4315
rect 358 4251 474 4315
rect 674 4251 790 4315
rect 990 4251 1106 4315
rect 1306 4251 1422 4315
rect 1622 4251 1738 4315
rect 1938 4251 2054 4315
rect 2254 4251 2370 4315
rect -3908 4126 -3792 4190
rect -3592 4126 -3476 4190
rect -3276 4126 -3160 4190
rect -2960 4126 -2844 4190
rect -2644 4126 -2528 4190
rect -2328 4126 -2212 4190
rect -2012 4126 -1896 4190
rect -1696 4126 -1580 4190
rect -1380 4126 -1264 4190
rect -1064 4126 -948 4190
rect -748 4126 -632 4190
rect -432 4126 -316 4190
rect -116 4126 0 4190
rect 200 4126 316 4190
rect 516 4126 632 4190
rect 832 4126 948 4190
rect 1148 4126 1264 4190
rect 1464 4126 1580 4190
rect 1780 4126 1896 4190
rect 2096 4126 2212 4190
rect -4118 3929 2350 3941
rect -4118 3889 2350 3929
rect -4118 3881 2350 3889
rect -4066 3631 -3950 3695
rect -3750 3631 -3634 3695
rect -3434 3631 -3318 3695
rect -3118 3631 -3002 3695
rect -2802 3631 -2686 3695
rect -2486 3631 -2370 3695
rect -2170 3631 -2054 3695
rect -1854 3631 -1738 3695
rect -1538 3631 -1422 3695
rect -1222 3631 -1106 3695
rect -906 3631 -790 3695
rect -590 3631 -474 3695
rect -274 3631 -158 3695
rect 42 3631 158 3695
rect 358 3631 474 3695
rect 674 3631 790 3695
rect 990 3631 1106 3695
rect 1306 3631 1422 3695
rect 1622 3631 1738 3695
rect 1938 3631 2054 3695
rect 2254 3631 2370 3695
rect -3908 3506 -3792 3570
rect -3592 3506 -3476 3570
rect -3276 3506 -3160 3570
rect -2960 3506 -2844 3570
rect -2644 3506 -2528 3570
rect -2328 3506 -2212 3570
rect -2012 3506 -1896 3570
rect -1696 3506 -1580 3570
rect -1380 3506 -1264 3570
rect -1064 3506 -948 3570
rect -748 3506 -632 3570
rect -432 3506 -316 3570
rect -116 3506 0 3570
rect 200 3506 316 3570
rect 516 3506 632 3570
rect 832 3506 948 3570
rect 1148 3506 1264 3570
rect 1464 3506 1580 3570
rect 1780 3506 1896 3570
rect 2096 3506 2212 3570
rect -4066 3196 -3950 3260
rect -3750 3196 -3634 3260
rect -3434 3196 -3318 3260
rect -3118 3196 -3002 3260
rect -2802 3196 -2686 3260
rect -2486 3196 -2370 3260
rect -2170 3196 -2054 3260
rect -1854 3196 -1738 3260
rect -1538 3196 -1422 3260
rect -1222 3196 -1106 3260
rect -906 3196 -790 3260
rect -590 3196 -474 3260
rect -274 3196 -158 3260
rect 42 3196 158 3260
rect 358 3196 474 3260
rect 674 3196 790 3260
rect 990 3196 1106 3260
rect 1306 3196 1422 3260
rect 1622 3196 1738 3260
rect 1938 3196 2054 3260
rect 2254 3196 2370 3260
rect -3908 3071 -3792 3135
rect -3592 3071 -3476 3135
rect -3276 3071 -3160 3135
rect -2960 3071 -2844 3135
rect -2644 3071 -2528 3135
rect -2328 3071 -2212 3135
rect -2012 3071 -1896 3135
rect -1696 3071 -1580 3135
rect -1380 3071 -1264 3135
rect -1064 3071 -948 3135
rect -748 3071 -632 3135
rect -432 3071 -316 3135
rect -116 3071 0 3135
rect 200 3071 316 3135
rect 516 3071 632 3135
rect 832 3071 948 3135
rect 1148 3071 1264 3135
rect 1464 3071 1580 3135
rect 1780 3071 1896 3135
rect 2096 3071 2212 3135
rect -4066 2761 -3950 2825
rect -3750 2761 -3634 2825
rect -3434 2761 -3318 2825
rect -3118 2761 -3002 2825
rect -2802 2761 -2686 2825
rect -2486 2761 -2370 2825
rect -2170 2761 -2054 2825
rect -1854 2761 -1738 2825
rect -1538 2761 -1422 2825
rect -1222 2761 -1106 2825
rect -906 2761 -790 2825
rect -590 2761 -474 2825
rect -274 2761 -158 2825
rect 42 2761 158 2825
rect 358 2761 474 2825
rect 674 2761 790 2825
rect 990 2761 1106 2825
rect 1306 2761 1422 2825
rect 1622 2761 1738 2825
rect 1938 2761 2054 2825
rect 2254 2761 2370 2825
rect -3908 2636 -3792 2700
rect -3592 2636 -3476 2700
rect -3276 2636 -3160 2700
rect -2960 2636 -2844 2700
rect -2644 2636 -2528 2700
rect -2328 2636 -2212 2700
rect -2012 2636 -1896 2700
rect -1696 2636 -1580 2700
rect -1380 2636 -1264 2700
rect -1064 2636 -948 2700
rect -748 2636 -632 2700
rect -432 2636 -316 2700
rect -116 2636 0 2700
rect 200 2636 316 2700
rect 516 2636 632 2700
rect 832 2636 948 2700
rect 1148 2636 1264 2700
rect 1464 2636 1580 2700
rect 1780 2636 1896 2700
rect 2096 2636 2212 2700
rect -4066 2326 -3950 2390
rect -3750 2326 -3634 2390
rect -3434 2326 -3318 2390
rect -3118 2326 -3002 2390
rect -2802 2326 -2686 2390
rect -2486 2326 -2370 2390
rect -2170 2326 -2054 2390
rect -1854 2326 -1738 2390
rect -1538 2326 -1422 2390
rect -1222 2326 -1106 2390
rect -906 2326 -790 2390
rect -590 2326 -474 2390
rect -274 2326 -158 2390
rect 42 2326 158 2390
rect 358 2326 474 2390
rect 674 2326 790 2390
rect 990 2326 1106 2390
rect 1306 2326 1422 2390
rect 1622 2326 1738 2390
rect 1938 2326 2054 2390
rect 2254 2326 2370 2390
rect -3908 2201 -3792 2265
rect -3592 2201 -3476 2265
rect -3276 2201 -3160 2265
rect -2960 2201 -2844 2265
rect -2644 2201 -2528 2265
rect -2328 2201 -2212 2265
rect -2012 2201 -1896 2265
rect -1696 2201 -1580 2265
rect -1380 2201 -1264 2265
rect -1064 2201 -948 2265
rect -748 2201 -632 2265
rect -432 2201 -316 2265
rect -116 2201 0 2265
rect 200 2201 316 2265
rect 516 2201 632 2265
rect 832 2201 948 2265
rect 1148 2201 1264 2265
rect 1464 2201 1580 2265
rect 1780 2201 1896 2265
rect 2096 2201 2212 2265
rect -4066 1891 -3950 1955
rect -3750 1891 -3634 1955
rect -3434 1891 -3318 1955
rect -3118 1891 -3002 1955
rect -2802 1891 -2686 1955
rect -2486 1891 -2370 1955
rect -2170 1891 -2054 1955
rect -1854 1891 -1738 1955
rect -1538 1891 -1422 1955
rect -1222 1891 -1106 1955
rect -906 1891 -790 1955
rect -590 1891 -474 1955
rect -274 1891 -158 1955
rect 42 1891 158 1955
rect 358 1891 474 1955
rect 674 1891 790 1955
rect 990 1891 1106 1955
rect 1306 1891 1422 1955
rect 1622 1891 1738 1955
rect 1938 1891 2054 1955
rect 2254 1891 2370 1955
rect -3908 1766 -3792 1830
rect -3592 1766 -3476 1830
rect -3276 1766 -3160 1830
rect -2960 1766 -2844 1830
rect -2644 1766 -2528 1830
rect -2328 1766 -2212 1830
rect -2012 1766 -1896 1830
rect -1696 1766 -1580 1830
rect -1380 1766 -1264 1830
rect -1064 1766 -948 1830
rect -748 1766 -632 1830
rect -432 1766 -316 1830
rect -116 1766 0 1830
rect 200 1766 316 1830
rect 516 1766 632 1830
rect 832 1766 948 1830
rect 1148 1766 1264 1830
rect 1464 1766 1580 1830
rect 1780 1766 1896 1830
rect 2096 1766 2212 1830
rect -4349 1120 -4156 1182
rect -4064 1190 -3828 1431
rect -4126 819 -3826 1019
rect -4994 468 -4930 578
rect -4994 -14 -4944 468
rect -4944 -14 -4930 468
rect -4680 -10 -4620 572
rect -4126 489 -3826 689
rect 2534 1506 2683 6106
rect -3185 1391 1307 1426
rect -3185 1236 1307 1391
rect -3185 1196 1307 1236
rect -3438 436 -3269 491
rect -2531 436 -2110 491
rect -3222 227 -3081 279
rect -4373 -308 -4134 2
rect -4882 -438 -4728 -348
rect -3829 22 -3774 167
rect -3892 -469 -3713 -408
rect -3214 -250 -3162 -69
rect -1356 434 -947 489
rect -2789 323 -2648 375
rect -2776 -250 -2724 -69
rect -1921 227 -1780 279
rect -2284 28 -2192 80
rect -2178 -247 -2126 -66
rect -1907 -248 -1855 -67
rect -1489 323 -1348 375
rect -1478 -247 -1426 -66
rect -611 648 -520 836
rect -657 323 -470 375
rect -981 28 -889 80
rect -26 646 65 834
rect -79 227 108 279
rect 396 646 487 834
rect 716 649 807 837
rect 986 659 1072 822
rect -874 -247 -822 -66
rect -713 -469 -559 -408
rect 250 -254 317 -85
rect 408 -234 475 -65
rect 569 -252 636 -83
rect 725 -234 792 -65
rect 887 -251 954 -82
rect 1035 -255 1107 -78
rect 1725 434 1966 489
rect 2127 1193 2347 1432
rect 1589 122 1726 174
rect 1320 -249 1387 -80
rect 1458 -324 1529 70
rect 2534 681 2683 1015
rect 2453 381 2683 616
rect 2453 -109 2683 126
rect -3681 -645 2244 -555
rect -4066 -942 -3950 -878
rect -3750 -942 -3634 -878
rect -3434 -942 -3318 -878
rect -3118 -942 -3002 -878
rect -2802 -942 -2686 -878
rect -2486 -942 -2370 -878
rect -2170 -942 -2054 -878
rect -1854 -942 -1738 -878
rect -1538 -942 -1422 -878
rect -1222 -942 -1106 -878
rect -906 -942 -790 -878
rect -590 -942 -474 -878
rect -274 -942 -158 -878
rect 42 -942 158 -878
rect 358 -942 474 -878
rect 674 -942 790 -878
rect 990 -942 1106 -878
rect 1306 -942 1422 -878
rect 1622 -942 1738 -878
rect 1938 -942 2054 -878
rect 2254 -942 2370 -878
rect -3908 -1067 -3792 -1003
rect -3592 -1067 -3476 -1003
rect -3276 -1067 -3160 -1003
rect -2960 -1067 -2844 -1003
rect -2644 -1067 -2528 -1003
rect -2328 -1067 -2212 -1003
rect -2012 -1067 -1896 -1003
rect -1696 -1067 -1580 -1003
rect -1380 -1067 -1264 -1003
rect -1064 -1067 -948 -1003
rect -748 -1067 -632 -1003
rect -432 -1067 -316 -1003
rect -116 -1067 0 -1003
rect 200 -1067 316 -1003
rect 516 -1067 632 -1003
rect 832 -1067 948 -1003
rect 1148 -1067 1264 -1003
rect 1464 -1067 1580 -1003
rect 1780 -1067 1896 -1003
rect 2096 -1067 2212 -1003
rect -4066 -1360 -3950 -1296
rect -3750 -1360 -3634 -1296
rect -3434 -1360 -3318 -1296
rect -3118 -1360 -3002 -1296
rect -2802 -1360 -2686 -1296
rect -2486 -1360 -2370 -1296
rect -2170 -1360 -2054 -1296
rect -1854 -1360 -1738 -1296
rect -1538 -1360 -1422 -1296
rect -1222 -1360 -1106 -1296
rect -906 -1360 -790 -1296
rect -590 -1360 -474 -1296
rect -274 -1360 -158 -1296
rect 42 -1360 158 -1296
rect 358 -1360 474 -1296
rect 674 -1360 790 -1296
rect 990 -1360 1106 -1296
rect 1306 -1360 1422 -1296
rect 1622 -1360 1738 -1296
rect 1938 -1360 2054 -1296
rect 2254 -1360 2370 -1296
rect -3908 -1485 -3792 -1421
rect -3592 -1485 -3476 -1421
rect -3276 -1485 -3160 -1421
rect -2960 -1485 -2844 -1421
rect -2644 -1485 -2528 -1421
rect -2328 -1485 -2212 -1421
rect -2012 -1485 -1896 -1421
rect -1696 -1485 -1580 -1421
rect -1380 -1485 -1264 -1421
rect -1064 -1485 -948 -1421
rect -748 -1485 -632 -1421
rect -432 -1485 -316 -1421
rect -116 -1485 0 -1421
rect 200 -1485 316 -1421
rect 516 -1485 632 -1421
rect 832 -1485 948 -1421
rect 1148 -1485 1264 -1421
rect 1464 -1485 1580 -1421
rect 1780 -1485 1896 -1421
rect 2096 -1485 2212 -1421
rect -4066 -1778 -3950 -1714
rect -3750 -1778 -3634 -1714
rect -3434 -1778 -3318 -1714
rect -3118 -1778 -3002 -1714
rect -2802 -1778 -2686 -1714
rect -2486 -1778 -2370 -1714
rect -2170 -1778 -2054 -1714
rect -1854 -1778 -1738 -1714
rect -1538 -1778 -1422 -1714
rect -1222 -1778 -1106 -1714
rect -906 -1778 -790 -1714
rect -590 -1778 -474 -1714
rect -274 -1778 -158 -1714
rect 42 -1778 158 -1714
rect 358 -1778 474 -1714
rect 674 -1778 790 -1714
rect 990 -1778 1106 -1714
rect 1306 -1778 1422 -1714
rect 1622 -1778 1738 -1714
rect 1938 -1778 2054 -1714
rect 2254 -1778 2370 -1714
rect -3908 -1903 -3792 -1839
rect -3592 -1903 -3476 -1839
rect -3276 -1903 -3160 -1839
rect -2960 -1903 -2844 -1839
rect -2644 -1903 -2528 -1839
rect -2328 -1903 -2212 -1839
rect -2012 -1903 -1896 -1839
rect -1696 -1903 -1580 -1839
rect -1380 -1903 -1264 -1839
rect -1064 -1903 -948 -1839
rect -748 -1903 -632 -1839
rect -432 -1903 -316 -1839
rect -116 -1903 0 -1839
rect 200 -1903 316 -1839
rect 516 -1903 632 -1839
rect 832 -1903 948 -1839
rect 1148 -1903 1264 -1839
rect 1464 -1903 1580 -1839
rect 1780 -1903 1896 -1839
rect 2096 -1903 2212 -1839
rect -4382 -2460 -4133 -2110
rect 1627 -3441 2200 -3267
rect 2629 -3231 2699 -3220
rect 2629 -3481 2685 -3231
rect 2685 -3481 2699 -3231
rect 2629 -3491 2699 -3481
<< metal2 >>
rect -4362 6488 2685 6535
rect -4362 6347 -4332 6488
rect 2644 6347 2685 6488
rect -4362 6313 2685 6347
rect -4362 5931 -4140 6313
rect -4081 6106 2683 6130
rect -4081 6055 2534 6106
rect -4081 5991 -4066 6055
rect -3950 5991 -3750 6055
rect -3634 5991 -3434 6055
rect -3318 5991 -3118 6055
rect -3002 5991 -2802 6055
rect -2686 5991 -2486 6055
rect -2370 5991 -2170 6055
rect -2054 5991 -1854 6055
rect -1738 5991 -1538 6055
rect -1422 5991 -1222 6055
rect -1106 5991 -906 6055
rect -790 5991 -590 6055
rect -474 5991 -274 6055
rect -158 5991 42 6055
rect 158 5991 358 6055
rect 474 5991 674 6055
rect 790 5991 990 6055
rect 1106 5991 1306 6055
rect 1422 5991 1622 6055
rect 1738 5991 1938 6055
rect 2054 5991 2254 6055
rect 2370 5991 2534 6055
rect -4362 5930 -4081 5931
rect -4362 5866 -3908 5930
rect -3792 5866 -3592 5930
rect -3476 5866 -3276 5930
rect -3160 5866 -2960 5930
rect -2844 5866 -2644 5930
rect -2528 5866 -2328 5930
rect -2212 5866 -2012 5930
rect -1896 5866 -1696 5930
rect -1580 5866 -1380 5930
rect -1264 5866 -1064 5930
rect -948 5866 -748 5930
rect -632 5866 -432 5930
rect -316 5866 -116 5930
rect 0 5866 200 5930
rect 316 5866 516 5930
rect 632 5866 832 5930
rect 948 5866 1148 5930
rect 1264 5866 1464 5930
rect 1580 5866 1780 5930
rect 1896 5866 2096 5930
rect 2212 5866 2399 5930
rect -4362 5792 2399 5866
rect -4362 5490 -4140 5792
rect -4081 5791 2399 5792
rect 2453 5690 2534 5991
rect -4081 5615 2534 5690
rect -4081 5551 -4066 5615
rect -3950 5551 -3750 5615
rect -3634 5551 -3434 5615
rect -3318 5551 -3118 5615
rect -3002 5551 -2802 5615
rect -2686 5551 -2486 5615
rect -2370 5551 -2170 5615
rect -2054 5551 -1854 5615
rect -1738 5551 -1538 5615
rect -1422 5551 -1222 5615
rect -1106 5551 -906 5615
rect -790 5551 -590 5615
rect -474 5551 -274 5615
rect -158 5551 42 5615
rect 158 5551 358 5615
rect 474 5551 674 5615
rect 790 5551 990 5615
rect 1106 5551 1306 5615
rect 1422 5551 1622 5615
rect 1738 5551 1938 5615
rect 2054 5551 2254 5615
rect 2370 5551 2534 5615
rect -4362 5426 -3908 5490
rect -3792 5426 -3592 5490
rect -3476 5426 -3276 5490
rect -3160 5426 -2960 5490
rect -2844 5426 -2644 5490
rect -2528 5426 -2328 5490
rect -2212 5426 -2012 5490
rect -1896 5426 -1696 5490
rect -1580 5426 -1380 5490
rect -1264 5426 -1064 5490
rect -948 5426 -748 5490
rect -632 5426 -432 5490
rect -316 5426 -116 5490
rect 0 5426 200 5490
rect 316 5426 516 5490
rect 632 5426 832 5490
rect 948 5426 1148 5490
rect 1264 5426 1464 5490
rect 1580 5426 1780 5490
rect 1896 5426 2096 5490
rect 2212 5426 2399 5490
rect -4362 5351 2399 5426
rect -4362 5050 -4140 5351
rect 2453 5250 2534 5551
rect -4081 5175 2534 5250
rect -4081 5111 -4066 5175
rect -3950 5111 -3750 5175
rect -3634 5111 -3434 5175
rect -3318 5111 -3118 5175
rect -3002 5111 -2802 5175
rect -2686 5111 -2486 5175
rect -2370 5111 -2170 5175
rect -2054 5111 -1854 5175
rect -1738 5111 -1538 5175
rect -1422 5111 -1222 5175
rect -1106 5111 -906 5175
rect -790 5111 -590 5175
rect -474 5111 -274 5175
rect -158 5111 42 5175
rect 158 5111 358 5175
rect 474 5111 674 5175
rect 790 5111 990 5175
rect 1106 5111 1306 5175
rect 1422 5111 1622 5175
rect 1738 5111 1938 5175
rect 2054 5111 2254 5175
rect 2370 5111 2534 5175
rect -4362 4986 -3908 5050
rect -3792 4986 -3592 5050
rect -3476 4986 -3276 5050
rect -3160 4986 -2960 5050
rect -2844 4986 -2644 5050
rect -2528 4986 -2328 5050
rect -2212 4986 -2012 5050
rect -1896 4986 -1696 5050
rect -1580 4986 -1380 5050
rect -1264 4986 -1064 5050
rect -948 4986 -748 5050
rect -632 4986 -432 5050
rect -316 4986 -116 5050
rect 0 4986 200 5050
rect 316 4986 516 5050
rect 632 4986 832 5050
rect 948 4986 1148 5050
rect 1264 4986 1464 5050
rect 1580 4986 1780 5050
rect 1896 4986 2096 5050
rect 2212 4986 2399 5050
rect -4362 4911 2399 4986
rect -4362 4615 -4140 4911
rect 2453 4815 2534 5111
rect -4081 4740 2534 4815
rect -4081 4676 -4066 4740
rect -3950 4676 -3750 4740
rect -3634 4676 -3434 4740
rect -3318 4676 -3118 4740
rect -3002 4676 -2802 4740
rect -2686 4676 -2486 4740
rect -2370 4676 -2170 4740
rect -2054 4676 -1854 4740
rect -1738 4676 -1538 4740
rect -1422 4676 -1222 4740
rect -1106 4676 -906 4740
rect -790 4676 -590 4740
rect -474 4676 -274 4740
rect -158 4676 42 4740
rect 158 4676 358 4740
rect 474 4676 674 4740
rect 790 4676 990 4740
rect 1106 4676 1306 4740
rect 1422 4676 1622 4740
rect 1738 4676 1938 4740
rect 2054 4676 2254 4740
rect 2370 4676 2534 4740
rect -4362 4551 -3908 4615
rect -3792 4551 -3592 4615
rect -3476 4551 -3276 4615
rect -3160 4551 -2960 4615
rect -2844 4551 -2644 4615
rect -2528 4551 -2328 4615
rect -2212 4551 -2012 4615
rect -1896 4551 -1696 4615
rect -1580 4551 -1380 4615
rect -1264 4551 -1064 4615
rect -948 4551 -748 4615
rect -632 4551 -432 4615
rect -316 4551 -116 4615
rect 0 4551 200 4615
rect 316 4551 516 4615
rect 632 4551 832 4615
rect 948 4551 1148 4615
rect 1264 4551 1464 4615
rect 1580 4551 1780 4615
rect 1896 4551 2096 4615
rect 2212 4551 2399 4615
rect -4362 4476 2399 4551
rect -4362 4190 -4140 4476
rect 2453 4390 2534 4676
rect -4081 4315 2534 4390
rect -4081 4251 -4066 4315
rect -3950 4251 -3750 4315
rect -3634 4251 -3434 4315
rect -3318 4251 -3118 4315
rect -3002 4251 -2802 4315
rect -2686 4251 -2486 4315
rect -2370 4251 -2170 4315
rect -2054 4251 -1854 4315
rect -1738 4251 -1538 4315
rect -1422 4251 -1222 4315
rect -1106 4251 -906 4315
rect -790 4251 -590 4315
rect -474 4251 -274 4315
rect -158 4251 42 4315
rect 158 4251 358 4315
rect 474 4251 674 4315
rect 790 4251 990 4315
rect 1106 4251 1306 4315
rect 1422 4251 1622 4315
rect 1738 4251 1938 4315
rect 2054 4251 2254 4315
rect 2370 4251 2534 4315
rect -4362 4126 -3908 4190
rect -3792 4126 -3592 4190
rect -3476 4126 -3276 4190
rect -3160 4126 -2960 4190
rect -2844 4126 -2644 4190
rect -2528 4126 -2328 4190
rect -2212 4126 -2012 4190
rect -1896 4126 -1696 4190
rect -1580 4126 -1380 4190
rect -1264 4126 -1064 4190
rect -948 4126 -748 4190
rect -632 4126 -432 4190
rect -316 4126 -116 4190
rect 0 4126 200 4190
rect 316 4126 516 4190
rect 632 4126 832 4190
rect 948 4126 1148 4190
rect 1264 4126 1464 4190
rect 1580 4126 1780 4190
rect 1896 4126 2096 4190
rect 2212 4126 2399 4190
rect -4362 4051 2399 4126
rect -4362 3941 -4140 4051
rect 2453 4002 2534 4251
rect 2470 3974 2534 4002
rect -4362 3881 -4118 3941
rect 2350 3881 2376 3941
rect -4362 3570 -4140 3881
rect 2453 3770 2534 3974
rect -4081 3695 2534 3770
rect -4081 3631 -4066 3695
rect -3950 3631 -3750 3695
rect -3634 3631 -3434 3695
rect -3318 3631 -3118 3695
rect -3002 3631 -2802 3695
rect -2686 3631 -2486 3695
rect -2370 3631 -2170 3695
rect -2054 3631 -1854 3695
rect -1738 3631 -1538 3695
rect -1422 3631 -1222 3695
rect -1106 3631 -906 3695
rect -790 3631 -590 3695
rect -474 3631 -274 3695
rect -158 3631 42 3695
rect 158 3631 358 3695
rect 474 3631 674 3695
rect 790 3631 990 3695
rect 1106 3631 1306 3695
rect 1422 3631 1622 3695
rect 1738 3631 1938 3695
rect 2054 3631 2254 3695
rect 2370 3631 2534 3695
rect -4362 3506 -3908 3570
rect -3792 3506 -3592 3570
rect -3476 3506 -3276 3570
rect -3160 3506 -2960 3570
rect -2844 3506 -2644 3570
rect -2528 3506 -2328 3570
rect -2212 3506 -2012 3570
rect -1896 3506 -1696 3570
rect -1580 3506 -1380 3570
rect -1264 3506 -1064 3570
rect -948 3506 -748 3570
rect -632 3506 -432 3570
rect -316 3506 -116 3570
rect 0 3506 200 3570
rect 316 3506 516 3570
rect 632 3506 832 3570
rect 948 3506 1148 3570
rect 1264 3506 1464 3570
rect 1580 3506 1780 3570
rect 1896 3506 2096 3570
rect 2212 3506 2399 3570
rect -4362 3431 2399 3506
rect -4362 3135 -4140 3431
rect 2453 3335 2534 3631
rect -4081 3260 2534 3335
rect -4081 3196 -4066 3260
rect -3950 3196 -3750 3260
rect -3634 3196 -3434 3260
rect -3318 3196 -3118 3260
rect -3002 3196 -2802 3260
rect -2686 3196 -2486 3260
rect -2370 3196 -2170 3260
rect -2054 3196 -1854 3260
rect -1738 3196 -1538 3260
rect -1422 3196 -1222 3260
rect -1106 3196 -906 3260
rect -790 3196 -590 3260
rect -474 3196 -274 3260
rect -158 3196 42 3260
rect 158 3196 358 3260
rect 474 3196 674 3260
rect 790 3196 990 3260
rect 1106 3196 1306 3260
rect 1422 3196 1622 3260
rect 1738 3196 1938 3260
rect 2054 3196 2254 3260
rect 2370 3196 2534 3260
rect -4362 3071 -3908 3135
rect -3792 3071 -3592 3135
rect -3476 3071 -3276 3135
rect -3160 3071 -2960 3135
rect -2844 3071 -2644 3135
rect -2528 3071 -2328 3135
rect -2212 3071 -2012 3135
rect -1896 3071 -1696 3135
rect -1580 3071 -1380 3135
rect -1264 3071 -1064 3135
rect -948 3071 -748 3135
rect -632 3071 -432 3135
rect -316 3071 -116 3135
rect 0 3071 200 3135
rect 316 3071 516 3135
rect 632 3071 832 3135
rect 948 3071 1148 3135
rect 1264 3071 1464 3135
rect 1580 3071 1780 3135
rect 1896 3071 2096 3135
rect 2212 3071 2399 3135
rect -4362 2996 2399 3071
rect -4362 2700 -4140 2996
rect 2453 2900 2534 3196
rect -4081 2825 2534 2900
rect -4081 2761 -4066 2825
rect -3950 2761 -3750 2825
rect -3634 2761 -3434 2825
rect -3318 2761 -3118 2825
rect -3002 2761 -2802 2825
rect -2686 2761 -2486 2825
rect -2370 2761 -2170 2825
rect -2054 2761 -1854 2825
rect -1738 2761 -1538 2825
rect -1422 2761 -1222 2825
rect -1106 2761 -906 2825
rect -790 2761 -590 2825
rect -474 2761 -274 2825
rect -158 2761 42 2825
rect 158 2761 358 2825
rect 474 2761 674 2825
rect 790 2761 990 2825
rect 1106 2761 1306 2825
rect 1422 2761 1622 2825
rect 1738 2761 1938 2825
rect 2054 2761 2254 2825
rect 2370 2761 2534 2825
rect -4362 2636 -3908 2700
rect -3792 2636 -3592 2700
rect -3476 2636 -3276 2700
rect -3160 2636 -2960 2700
rect -2844 2636 -2644 2700
rect -2528 2636 -2328 2700
rect -2212 2636 -2012 2700
rect -1896 2636 -1696 2700
rect -1580 2636 -1380 2700
rect -1264 2636 -1064 2700
rect -948 2636 -748 2700
rect -632 2636 -432 2700
rect -316 2636 -116 2700
rect 0 2636 200 2700
rect 316 2636 516 2700
rect 632 2636 832 2700
rect 948 2636 1148 2700
rect 1264 2636 1464 2700
rect 1580 2636 1780 2700
rect 1896 2636 2096 2700
rect 2212 2636 2399 2700
rect -4362 2561 2399 2636
rect -4362 2265 -4140 2561
rect 2453 2465 2534 2761
rect -4081 2390 2534 2465
rect -4081 2326 -4066 2390
rect -3950 2326 -3750 2390
rect -3634 2326 -3434 2390
rect -3318 2326 -3118 2390
rect -3002 2326 -2802 2390
rect -2686 2326 -2486 2390
rect -2370 2326 -2170 2390
rect -2054 2326 -1854 2390
rect -1738 2326 -1538 2390
rect -1422 2326 -1222 2390
rect -1106 2326 -906 2390
rect -790 2326 -590 2390
rect -474 2326 -274 2390
rect -158 2326 42 2390
rect 158 2326 358 2390
rect 474 2326 674 2390
rect 790 2326 990 2390
rect 1106 2326 1306 2390
rect 1422 2326 1622 2390
rect 1738 2326 1938 2390
rect 2054 2326 2254 2390
rect 2370 2326 2534 2390
rect -4362 2201 -3908 2265
rect -3792 2201 -3592 2265
rect -3476 2201 -3276 2265
rect -3160 2201 -2960 2265
rect -2844 2201 -2644 2265
rect -2528 2201 -2328 2265
rect -2212 2201 -2012 2265
rect -1896 2201 -1696 2265
rect -1580 2201 -1380 2265
rect -1264 2201 -1064 2265
rect -948 2201 -748 2265
rect -632 2201 -432 2265
rect -316 2201 -116 2265
rect 0 2201 200 2265
rect 316 2201 516 2265
rect 632 2201 832 2265
rect 948 2201 1148 2265
rect 1264 2201 1464 2265
rect 1580 2201 1780 2265
rect 1896 2201 2096 2265
rect 2212 2201 2399 2265
rect -4362 2126 2399 2201
rect -4362 1830 -4140 2126
rect 2453 2030 2534 2326
rect -4081 1955 2534 2030
rect -4081 1891 -4066 1955
rect -3950 1891 -3750 1955
rect -3634 1891 -3434 1955
rect -3318 1891 -3118 1955
rect -3002 1891 -2802 1955
rect -2686 1891 -2486 1955
rect -2370 1891 -2170 1955
rect -2054 1891 -1854 1955
rect -1738 1891 -1538 1955
rect -1422 1891 -1222 1955
rect -1106 1891 -906 1955
rect -790 1891 -590 1955
rect -474 1891 -274 1955
rect -158 1891 42 1955
rect 158 1891 358 1955
rect 474 1891 674 1955
rect 790 1891 990 1955
rect 1106 1891 1306 1955
rect 1422 1891 1622 1955
rect 1738 1891 1938 1955
rect 2054 1891 2254 1955
rect 2370 1891 2534 1955
rect -4362 1766 -3908 1830
rect -3792 1766 -3592 1830
rect -3476 1766 -3276 1830
rect -3160 1766 -2960 1830
rect -2844 1766 -2644 1830
rect -2528 1766 -2328 1830
rect -2212 1766 -2012 1830
rect -1896 1766 -1696 1830
rect -1580 1766 -1380 1830
rect -1264 1766 -1064 1830
rect -948 1766 -748 1830
rect -632 1766 -432 1830
rect -316 1766 -116 1830
rect 0 1766 200 1830
rect 316 1766 516 1830
rect 632 1766 832 1830
rect 948 1766 1148 1830
rect 1264 1766 1464 1830
rect 1580 1766 1780 1830
rect 1896 1766 2096 1830
rect 2212 1766 2399 1830
rect -4362 1691 2399 1766
rect -4362 1445 -4140 1691
rect 2453 1506 2534 1891
rect -4362 1432 2363 1445
rect -4362 1431 2127 1432
rect -4362 1190 -4064 1431
rect -3828 1426 2127 1431
rect -3828 1196 -3185 1426
rect 1307 1196 2127 1426
rect -3828 1193 2127 1196
rect 2347 1193 2363 1432
rect -3828 1190 2363 1193
rect -4362 1182 2363 1190
rect -4362 1120 -4349 1182
rect -4156 1177 2363 1182
rect -4156 1120 -4140 1177
rect -4362 1106 -4140 1120
rect -5034 588 -4932 862
rect -5034 578 -4930 588
rect -5034 -14 -4994 578
rect -5034 -24 -4930 -14
rect -4680 572 -4542 862
rect -4144 819 -4126 1019
rect -3826 874 -3808 1019
rect -3826 819 -3513 874
rect -4620 -10 -4542 572
rect -4144 489 -4126 689
rect -3826 277 -3762 689
rect -3568 373 -3513 819
rect -783 837 821 847
rect -783 836 716 837
rect -783 648 -611 836
rect -520 834 716 836
rect -520 648 -26 834
rect -783 646 -26 648
rect 65 646 396 834
rect 487 649 716 834
rect 807 649 821 837
rect 977 822 1082 1177
rect 977 659 986 822
rect 1072 659 1082 822
rect 977 652 1082 659
rect 2453 1015 2683 1506
rect 2453 681 2534 1015
rect 487 646 821 649
rect -783 637 821 646
rect 2453 633 2683 681
rect 2453 616 2699 633
rect -3445 436 -3438 491
rect -3269 436 -2531 491
rect -2110 436 -2097 491
rect -1377 434 -1356 489
rect -947 434 1725 489
rect 1966 434 1975 489
rect 2683 381 2699 616
rect -2795 373 -2789 375
rect -3568 323 -2789 373
rect -2648 373 -2642 375
rect -1495 373 -1489 375
rect -2648 323 -1489 373
rect -1348 373 -1342 375
rect -665 373 -657 375
rect -1348 323 -657 373
rect -470 323 -461 375
rect -3228 277 -3222 279
rect -3826 227 -3222 277
rect -3081 277 -3075 279
rect -1927 277 -1921 279
rect -3081 227 -1921 277
rect -1780 277 -1774 279
rect -89 277 -79 279
rect -1780 227 -79 277
rect 108 227 118 279
rect -89 224 118 227
rect -3829 167 1589 174
rect -5034 -348 -4932 -24
rect -4882 -348 -4728 -338
rect -4680 -348 -4542 -10
rect -4392 2 -4121 44
rect -3774 132 1589 167
rect 1583 122 1589 132
rect 1726 122 1732 174
rect 2453 126 2699 381
rect -2293 28 -2284 80
rect -2192 70 -2186 80
rect -987 70 -981 80
rect -2192 28 -981 70
rect -889 70 -883 80
rect 1458 70 1529 78
rect -889 28 1458 70
rect -3829 15 -3774 22
rect -4392 -308 -4373 2
rect -4134 -308 -4121 2
rect -3221 -66 -2118 -60
rect -3221 -69 -2178 -66
rect -3221 -250 -3214 -69
rect -3162 -250 -2776 -69
rect -2724 -247 -2178 -69
rect -2126 -247 -2118 -66
rect -2724 -250 -2118 -247
rect -3221 -256 -2118 -250
rect -1916 -66 -816 -60
rect -1916 -67 -1478 -66
rect -1916 -248 -1907 -67
rect -1855 -247 -1478 -67
rect -1426 -247 -874 -66
rect -822 -247 -816 -66
rect 397 -65 485 28
rect -1855 -248 -816 -247
rect -1916 -256 -816 -248
rect 239 -85 326 -79
rect 239 -254 250 -85
rect 317 -254 326 -85
rect 397 -234 408 -65
rect 475 -234 485 -65
rect 717 -65 805 28
rect 397 -243 485 -234
rect 560 -83 647 -72
rect -4392 -348 -4121 -308
rect -5034 -396 -4882 -348
rect -5032 -438 -4882 -396
rect -4728 -438 -4121 -348
rect -5032 -531 -4121 -438
rect -3909 -469 -3892 -408
rect -3713 -469 -713 -408
rect -559 -469 -551 -408
rect 239 -531 326 -254
rect 560 -252 569 -83
rect 636 -252 647 -83
rect 717 -234 725 -65
rect 792 -234 805 -65
rect 717 -243 805 -234
rect 879 -82 966 -72
rect 560 -531 647 -252
rect 879 -251 887 -82
rect 954 -251 966 -82
rect 879 -531 966 -251
rect 1028 -78 1115 28
rect 1028 -255 1035 -78
rect 1107 -255 1115 -78
rect 1028 -330 1115 -255
rect 1312 -80 1399 -73
rect 1312 -249 1320 -80
rect 1387 -249 1399 -80
rect 1312 -531 1399 -249
rect 1458 -337 1529 -324
rect 2683 -109 2699 126
rect -5032 -555 2271 -531
rect -5032 -580 -3681 -555
rect -4680 -582 -4542 -580
rect -4392 -645 -3681 -580
rect 2244 -645 2271 -555
rect -4392 -685 2271 -645
rect -4392 -1003 -4121 -685
rect 2453 -803 2699 -109
rect -4092 -878 2699 -803
rect -4092 -942 -4066 -878
rect -3950 -942 -3750 -878
rect -3634 -942 -3434 -878
rect -3318 -942 -3118 -878
rect -3002 -942 -2802 -878
rect -2686 -942 -2486 -878
rect -2370 -942 -2170 -878
rect -2054 -942 -1854 -878
rect -1738 -942 -1538 -878
rect -1422 -942 -1222 -878
rect -1106 -942 -906 -878
rect -790 -942 -590 -878
rect -474 -942 -274 -878
rect -158 -942 42 -878
rect 158 -942 358 -878
rect 474 -942 674 -878
rect 790 -942 990 -878
rect 1106 -942 1306 -878
rect 1422 -942 1622 -878
rect 1738 -942 1938 -878
rect 2054 -942 2254 -878
rect 2370 -942 2699 -878
rect -4393 -1067 -3908 -1003
rect -3792 -1067 -3592 -1003
rect -3476 -1067 -3276 -1003
rect -3160 -1067 -2960 -1003
rect -2844 -1067 -2644 -1003
rect -2528 -1067 -2328 -1003
rect -2212 -1067 -2012 -1003
rect -1896 -1067 -1696 -1003
rect -1580 -1067 -1380 -1003
rect -1264 -1067 -1064 -1003
rect -948 -1067 -748 -1003
rect -632 -1067 -432 -1003
rect -316 -1067 -116 -1003
rect 0 -1067 200 -1003
rect 316 -1067 516 -1003
rect 632 -1067 832 -1003
rect 948 -1067 1148 -1003
rect 1264 -1067 1464 -1003
rect 1580 -1067 1780 -1003
rect 1896 -1067 2096 -1003
rect 2212 -1067 2383 -1003
rect -4393 -1142 2383 -1067
rect -4392 -1421 -4121 -1142
rect 2437 -1221 2699 -942
rect -4081 -1296 2699 -1221
rect -4081 -1360 -4066 -1296
rect -3950 -1360 -3750 -1296
rect -3634 -1360 -3434 -1296
rect -3318 -1360 -3118 -1296
rect -3002 -1360 -2802 -1296
rect -2686 -1360 -2486 -1296
rect -2370 -1360 -2170 -1296
rect -2054 -1360 -1854 -1296
rect -1738 -1360 -1538 -1296
rect -1422 -1360 -1222 -1296
rect -1106 -1360 -906 -1296
rect -790 -1360 -590 -1296
rect -474 -1360 -274 -1296
rect -158 -1360 42 -1296
rect 158 -1360 358 -1296
rect 474 -1360 674 -1296
rect 790 -1360 990 -1296
rect 1106 -1360 1306 -1296
rect 1422 -1360 1622 -1296
rect 1738 -1360 1938 -1296
rect 2054 -1360 2254 -1296
rect 2370 -1360 2699 -1296
rect -4392 -1485 -3908 -1421
rect -3792 -1485 -3592 -1421
rect -3476 -1485 -3276 -1421
rect -3160 -1485 -2960 -1421
rect -2844 -1485 -2644 -1421
rect -2528 -1485 -2328 -1421
rect -2212 -1485 -2012 -1421
rect -1896 -1485 -1696 -1421
rect -1580 -1485 -1380 -1421
rect -1264 -1485 -1064 -1421
rect -948 -1485 -748 -1421
rect -632 -1485 -432 -1421
rect -316 -1485 -116 -1421
rect 0 -1485 200 -1421
rect 316 -1485 516 -1421
rect 632 -1485 832 -1421
rect 948 -1485 1148 -1421
rect 1264 -1485 1464 -1421
rect 1580 -1485 1780 -1421
rect 1896 -1485 2096 -1421
rect 2212 -1485 2383 -1421
rect -4392 -1560 2383 -1485
rect -4392 -1839 -4121 -1560
rect 2437 -1639 2699 -1360
rect -4081 -1714 2699 -1639
rect -4081 -1778 -4066 -1714
rect -3950 -1778 -3750 -1714
rect -3634 -1778 -3434 -1714
rect -3318 -1778 -3118 -1714
rect -3002 -1778 -2802 -1714
rect -2686 -1778 -2486 -1714
rect -2370 -1778 -2170 -1714
rect -2054 -1778 -1854 -1714
rect -1738 -1778 -1538 -1714
rect -1422 -1778 -1222 -1714
rect -1106 -1778 -906 -1714
rect -790 -1778 -590 -1714
rect -474 -1778 -274 -1714
rect -158 -1778 42 -1714
rect 158 -1778 358 -1714
rect 474 -1778 674 -1714
rect 790 -1778 990 -1714
rect 1106 -1778 1306 -1714
rect 1422 -1778 1622 -1714
rect 1738 -1778 1938 -1714
rect 2054 -1778 2254 -1714
rect 2370 -1778 2699 -1714
rect -4392 -1903 -3908 -1839
rect -3792 -1903 -3592 -1839
rect -3476 -1903 -3276 -1839
rect -3160 -1903 -2960 -1839
rect -2844 -1903 -2644 -1839
rect -2528 -1903 -2328 -1839
rect -2212 -1903 -2012 -1839
rect -1896 -1903 -1696 -1839
rect -1580 -1903 -1380 -1839
rect -1264 -1903 -1064 -1839
rect -948 -1903 -748 -1839
rect -632 -1903 -432 -1839
rect -316 -1903 -116 -1839
rect 0 -1903 200 -1839
rect 316 -1903 516 -1839
rect 632 -1903 832 -1839
rect 948 -1903 1148 -1839
rect 1264 -1903 1464 -1839
rect 1580 -1903 1780 -1839
rect 1896 -1903 2096 -1839
rect 2212 -1903 2383 -1839
rect -4392 -1978 2383 -1903
rect -4392 -2110 -4121 -1978
rect -4392 -2460 -4382 -2110
rect -4133 -2460 -4121 -2110
rect -4392 -2472 -4121 -2460
rect 1573 -3267 2629 -3220
rect 1573 -3441 1627 -3267
rect 2200 -3441 2629 -3267
rect 1573 -3491 2629 -3441
rect 2699 -3491 2705 -3220
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  M13 ~/Tesis/magic/buffer/paramcells
timestamp 1652924542
transform 1 0 1710 0 1 -157
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  M24
timestamp 1652924542
transform 1 0 1275 0 1 -157
box -278 -358 278 358
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_0 ~/Tesis/magic/buffer/paramcells
timestamp 1652928066
transform 1 0 -3804 0 1 -100
box -198 -198 198 198
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_1
timestamp 1652928066
transform 1 0 -3804 0 1 500
box -198 -198 198 198
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_2
timestamp 1652928066
transform 1 0 -3804 0 1 915
box -198 -198 198 198
use sky130_fd_pr__nfet_03v3_nvt_EJGQJV  sky130_fd_pr__nfet_03v3_nvt_EJGQJV_0 ~/Tesis/magic/buffer/paramcells
timestamp 1652924542
transform -1 0 -2671 0 1 -157
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_AQ2AJT  sky130_fd_pr__pfet_g5v0d10v5_AQ2AJT_0 ~/Tesis/magic/buffer/paramcells
timestamp 1652924542
transform 1 0 -849 0 1 5083
box -3389 -1269 3389 1269
use sky130_fd_pr__pfet_g5v0d10v5_AQ2AJT  sky130_fd_pr__pfet_g5v0d10v5_AQ2AJT_1
timestamp 1652924542
transform 1 0 -849 0 1 2735
box -3389 -1269 3389 1269
use sky130_fd_pr__res_xhigh_po_0p35_D7NTZ8  sky130_fd_pr__res_xhigh_po_0p35_D7NTZ8_0 ~/Tesis/magic/buffer/paramcells
timestamp 1652924542
transform 0 1 -890 -1 0 -2878
box -678 -3098 678 3098
use sky130_fd_pr__res_xhigh_po_0p35_HT39D6  sky130_fd_pr__res_xhigh_po_0p35_HT39D6_1 ~/Tesis/magic/buffer/paramcells
timestamp 1723585349
transform 1 0 -4807 0 1 259
box -201 -683 201 683
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM1
timestamp 1652924542
transform -1 0 -1803 0 1 -157
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM2
timestamp 1652924542
transform -1 0 -1369 0 1 -157
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM3 ~/Tesis/magic/buffer/paramcells
timestamp 1652924542
transform 1 0 -2319 0 1 704
box -387 -362 387 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM4
timestamp 1652924542
transform -1 0 -1151 0 1 704
box -387 -362 387 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM5
timestamp 1652924542
transform -1 0 -1735 0 1 704
box -387 -362 387 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM6
timestamp 1652924542
transform 1 0 -2903 0 1 704
box -387 -362 387 362
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM7
timestamp 1652924542
transform -1 0 -2237 0 1 -157
box -278 -358 278 358
use sky130_fd_pr__nfet_03v3_nvt_EJGQJV  XM8
timestamp 1652924542
transform -1 0 -3105 0 1 -157
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM9
timestamp 1652924542
transform -1 0 -935 0 1 -157
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_H7BQ24  XM10 ~/Tesis/magic/buffer/paramcells
timestamp 1723585349
transform 1 0 603 0 1 -158
box -515 -358 515 358
use sky130_fd_pr__nfet_g5v0d10v5_UC3VEF  XM22 ~/Tesis/magic/buffer/paramcells
timestamp 1652924542
transform 1 0 -865 0 1 -1392
box -3359 -776 3359 776
use sky130_fd_pr__pfet_g5v0d10v5_U6NWY6  XM25 ~/Tesis/magic/buffer/paramcells
timestamp 1652924542
transform 1 0 1106 0 1 704
box -308 -362 308 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM26
timestamp 1652924542
transform 1 0 601 0 1 704
box -387 -362 387 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM27
timestamp 1652924542
transform 1 0 17 0 1 704
box -387 -362 387 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM28
timestamp 1652924542
transform 1 0 -567 0 1 704
box -387 -362 387 362
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM29
timestamp 1652924542
transform -1 0 -501 0 1 -157
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM30
timestamp 1652924542
transform -1 0 -67 0 1 -157
box -278 -358 278 358
<< labels >>
flabel metal1 -4342 1201 -4142 1401 0 FreeSans 256 0 0 0 vdd
port 1 nsew
flabel metal1 2467 163 2667 363 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal2 -241 738 -241 738 0 FreeSans 320 0 0 0 vcomp
flabel metal2 -3529 -437 -3529 -437 0 FreeSans 320 0 0 0 ndrv
flabel metal2 1374 46 1374 46 0 FreeSans 320 0 0 0 nbias
flabel metal1 980 577 980 577 0 FreeSans 320 0 0 0 pbias
flabel metal2 -2456 -160 -2456 -160 0 FreeSans 320 0 0 0 vcomn2
flabel metal2 -1322 -168 -1322 -168 0 FreeSans 320 0 0 0 vcomn1
flabel metal1 -4361 164 -4161 364 0 FreeSans 320 0 0 0 ena
port 3 nsew
flabel metal2 1468 463 1468 463 0 FreeSans 320 0 0 0 pdrv1
flabel metal2 -3236 462 -3236 462 0 FreeSans 320 0 0 0 pdrv2
flabel metal1 -4361 489 -4161 689 0 FreeSans 256 0 0 0 inm
port 6 nsew
flabel metal1 -4361 819 -4161 1019 0 FreeSans 256 0 0 0 inp
port 5 nsew
flabel metal1 -4355 -529 -4155 -329 0 FreeSans 256 0 0 0 vss
port 4 nsew
<< end >>
