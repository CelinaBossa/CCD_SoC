magic
tech sky130A
magscale 1 2
timestamp 1723064828
<< nwell >>
rect -387 -397 387 397
<< mvpmos >>
rect -129 -100 -29 100
rect 29 -100 129 100
<< mvpdiff >>
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
<< mvpdiffc >>
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
<< mvnsubdiff >>
rect -321 319 321 331
rect -321 285 -213 319
rect 213 285 321 319
rect -321 273 321 285
rect -321 223 -263 273
rect -321 -223 -309 223
rect -275 -223 -263 223
rect 263 223 321 273
rect -321 -273 -263 -223
rect 263 -223 275 223
rect 309 -223 321 223
rect 263 -273 321 -223
rect -321 -285 321 -273
rect -321 -319 -213 -285
rect 213 -319 321 -285
rect -321 -331 321 -319
<< mvnsubdiffcont >>
rect -213 285 213 319
rect -309 -223 -275 223
rect 275 -223 309 223
rect -213 -319 213 -285
<< poly >>
rect -129 181 -29 197
rect -129 147 -113 181
rect -45 147 -29 181
rect -129 100 -29 147
rect 29 181 129 197
rect 29 147 45 181
rect 113 147 129 181
rect 29 100 129 147
rect -129 -147 -29 -100
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect -129 -197 -29 -181
rect 29 -147 129 -100
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 29 -197 129 -181
<< polycont >>
rect -113 147 -45 181
rect 45 147 113 181
rect -113 -181 -45 -147
rect 45 -181 113 -147
<< locali >>
rect -309 285 -213 319
rect 213 285 309 319
rect -309 223 -275 285
rect 275 223 309 285
rect -129 147 -113 181
rect -45 147 -29 181
rect 29 147 45 181
rect 113 147 129 181
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 113 -181 129 -147
rect -309 -285 -275 -223
rect 275 -285 309 -223
rect -309 -319 -213 -285
rect 213 -319 309 -285
<< viali >>
rect -113 147 -45 181
rect 45 147 113 181
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect -113 -181 -45 -147
rect 45 -181 113 -147
<< metal1 >>
rect -125 181 -33 187
rect -125 147 -113 181
rect -45 147 -33 181
rect -125 141 -33 147
rect 33 181 125 187
rect 33 147 45 181
rect 113 147 125 181
rect 33 141 125 147
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect -125 -147 -33 -141
rect -125 -181 -113 -147
rect -45 -181 -33 -147
rect -125 -187 -33 -181
rect 33 -147 125 -141
rect 33 -181 45 -147
rect 113 -181 125 -147
rect 33 -187 125 -181
<< properties >>
string FIXED_BBOX -292 -302 292 302
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
