magic
tech sky130A
magscale 1 2
timestamp 1723067318
<< locali >>
rect -30 553 30 610
rect -30 -610 30 -553
<< rlocali >>
rect -30 -553 30 553
<< properties >>
string gencell sky130_fd_pr__res_generic_l1
string library sky130
string parameters w 0.3 l 5.533 m 1 nx 1 wmin 0.17 lmin 0.17 rho 12.8 val 236.074 dummy 0 dw 0.0 term 0.0 snake 0 roverlap 0
<< end >>
