VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__opamp
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__opamp ;
  ORIGIN 31.350 24.580 ;
  SIZE 52.910 BY 62.500 ;
  PIN vdd
    ANTENNADIFFAREA 186.130493 ;
    PORT
      LAYER nwell ;
        RECT -22.735 7.330 14.085 33.205 ;
        RECT -22.735 -17.930 -21.160 7.330 ;
        RECT -16.450 1.710 7.070 5.330 ;
        RECT 12.510 -17.930 14.085 7.330 ;
        RECT -22.735 -19.505 14.085 -17.930 ;
      LAYER li1 ;
        RECT -22.305 31.200 13.655 32.775 ;
        RECT -22.305 19.645 -20.630 31.200 ;
        RECT -19.340 29.255 -19.170 30.295 ;
        RECT -17.760 29.255 -17.590 30.295 ;
        RECT -16.180 29.255 -16.010 30.295 ;
        RECT -14.600 29.255 -14.430 30.295 ;
        RECT -13.020 29.255 -12.850 30.295 ;
        RECT -11.440 29.255 -11.270 30.295 ;
        RECT -9.860 29.255 -9.690 30.295 ;
        RECT -8.280 29.255 -8.110 30.295 ;
        RECT -6.700 29.255 -6.530 30.295 ;
        RECT -5.120 29.255 -4.950 30.295 ;
        RECT -3.540 29.255 -3.370 30.295 ;
        RECT -1.960 29.255 -1.790 30.295 ;
        RECT -0.380 29.255 -0.210 30.295 ;
        RECT 1.200 29.255 1.370 30.295 ;
        RECT 2.780 29.255 2.950 30.295 ;
        RECT 4.360 29.255 4.530 30.295 ;
        RECT 5.940 29.255 6.110 30.295 ;
        RECT 7.520 29.255 7.690 30.295 ;
        RECT 9.100 29.255 9.270 30.295 ;
        RECT 10.680 29.255 10.850 30.295 ;
        RECT -19.340 27.075 -19.170 28.115 ;
        RECT -17.760 27.075 -17.590 28.115 ;
        RECT -16.180 27.075 -16.010 28.115 ;
        RECT -14.600 27.075 -14.430 28.115 ;
        RECT -13.020 27.075 -12.850 28.115 ;
        RECT -11.440 27.075 -11.270 28.115 ;
        RECT -9.860 27.075 -9.690 28.115 ;
        RECT -8.280 27.075 -8.110 28.115 ;
        RECT -6.700 27.075 -6.530 28.115 ;
        RECT -5.120 27.075 -4.950 28.115 ;
        RECT -3.540 27.075 -3.370 28.115 ;
        RECT -1.960 27.075 -1.790 28.115 ;
        RECT -0.380 27.075 -0.210 28.115 ;
        RECT 1.200 27.075 1.370 28.115 ;
        RECT 2.780 27.075 2.950 28.115 ;
        RECT 4.360 27.075 4.530 28.115 ;
        RECT 5.940 27.075 6.110 28.115 ;
        RECT 7.520 27.075 7.690 28.115 ;
        RECT 9.100 27.075 9.270 28.115 ;
        RECT 10.680 27.075 10.850 28.115 ;
        RECT -19.340 24.895 -19.170 25.935 ;
        RECT -17.760 24.895 -17.590 25.935 ;
        RECT -16.180 24.895 -16.010 25.935 ;
        RECT -14.600 24.895 -14.430 25.935 ;
        RECT -13.020 24.895 -12.850 25.935 ;
        RECT -11.440 24.895 -11.270 25.935 ;
        RECT -9.860 24.895 -9.690 25.935 ;
        RECT -8.280 24.895 -8.110 25.935 ;
        RECT -6.700 24.895 -6.530 25.935 ;
        RECT -5.120 24.895 -4.950 25.935 ;
        RECT -3.540 24.895 -3.370 25.935 ;
        RECT -1.960 24.895 -1.790 25.935 ;
        RECT -0.380 24.895 -0.210 25.935 ;
        RECT 1.200 24.895 1.370 25.935 ;
        RECT 2.780 24.895 2.950 25.935 ;
        RECT 4.360 24.895 4.530 25.935 ;
        RECT 5.940 24.895 6.110 25.935 ;
        RECT 7.520 24.895 7.690 25.935 ;
        RECT 9.100 24.895 9.270 25.935 ;
        RECT 10.680 24.895 10.850 25.935 ;
        RECT -19.340 22.715 -19.170 23.755 ;
        RECT -17.760 22.715 -17.590 23.755 ;
        RECT -16.180 22.715 -16.010 23.755 ;
        RECT -14.600 22.715 -14.430 23.755 ;
        RECT -13.020 22.715 -12.850 23.755 ;
        RECT -11.440 22.715 -11.270 23.755 ;
        RECT -9.860 22.715 -9.690 23.755 ;
        RECT -8.280 22.715 -8.110 23.755 ;
        RECT -6.700 22.715 -6.530 23.755 ;
        RECT -5.120 22.715 -4.950 23.755 ;
        RECT -3.540 22.715 -3.370 23.755 ;
        RECT -1.960 22.715 -1.790 23.755 ;
        RECT -0.380 22.715 -0.210 23.755 ;
        RECT 1.200 22.715 1.370 23.755 ;
        RECT 2.780 22.715 2.950 23.755 ;
        RECT 4.360 22.715 4.530 23.755 ;
        RECT 5.940 22.715 6.110 23.755 ;
        RECT 7.520 22.715 7.690 23.755 ;
        RECT 9.100 22.715 9.270 23.755 ;
        RECT 10.680 22.715 10.850 23.755 ;
        RECT -19.340 20.535 -19.170 21.575 ;
        RECT -17.760 20.535 -17.590 21.575 ;
        RECT -16.180 20.535 -16.010 21.575 ;
        RECT -14.600 20.535 -14.430 21.575 ;
        RECT -13.020 20.535 -12.850 21.575 ;
        RECT -11.440 20.535 -11.270 21.575 ;
        RECT -9.860 20.535 -9.690 21.575 ;
        RECT -8.280 20.535 -8.110 21.575 ;
        RECT -6.700 20.535 -6.530 21.575 ;
        RECT -5.120 20.535 -4.950 21.575 ;
        RECT -3.540 20.535 -3.370 21.575 ;
        RECT -1.960 20.535 -1.790 21.575 ;
        RECT -0.380 20.535 -0.210 21.575 ;
        RECT 1.200 20.535 1.370 21.575 ;
        RECT 2.780 20.535 2.950 21.575 ;
        RECT 4.360 20.535 4.530 21.575 ;
        RECT 5.940 20.535 6.110 21.575 ;
        RECT 7.520 20.535 7.690 21.575 ;
        RECT 9.100 20.535 9.270 21.575 ;
        RECT 10.680 20.535 10.850 21.575 ;
        RECT 12.140 19.645 13.655 31.200 ;
        RECT -22.305 19.445 13.655 19.645 ;
        RECT -22.305 7.890 -20.630 19.445 ;
        RECT -19.340 17.515 -19.170 18.555 ;
        RECT -17.760 17.515 -17.590 18.555 ;
        RECT -16.180 17.515 -16.010 18.555 ;
        RECT -14.600 17.515 -14.430 18.555 ;
        RECT -13.020 17.515 -12.850 18.555 ;
        RECT -11.440 17.515 -11.270 18.555 ;
        RECT -9.860 17.515 -9.690 18.555 ;
        RECT -8.280 17.515 -8.110 18.555 ;
        RECT -6.700 17.515 -6.530 18.555 ;
        RECT -5.120 17.515 -4.950 18.555 ;
        RECT -3.540 17.515 -3.370 18.555 ;
        RECT -1.960 17.515 -1.790 18.555 ;
        RECT -0.380 17.515 -0.210 18.555 ;
        RECT 1.200 17.515 1.370 18.555 ;
        RECT 2.780 17.515 2.950 18.555 ;
        RECT 4.360 17.515 4.530 18.555 ;
        RECT 5.940 17.515 6.110 18.555 ;
        RECT 7.520 17.515 7.690 18.555 ;
        RECT 9.100 17.515 9.270 18.555 ;
        RECT 10.680 17.515 10.850 18.555 ;
        RECT -19.340 15.335 -19.170 16.375 ;
        RECT -17.760 15.335 -17.590 16.375 ;
        RECT -16.180 15.335 -16.010 16.375 ;
        RECT -14.600 15.335 -14.430 16.375 ;
        RECT -13.020 15.335 -12.850 16.375 ;
        RECT -11.440 15.335 -11.270 16.375 ;
        RECT -9.860 15.335 -9.690 16.375 ;
        RECT -8.280 15.335 -8.110 16.375 ;
        RECT -6.700 15.335 -6.530 16.375 ;
        RECT -5.120 15.335 -4.950 16.375 ;
        RECT -3.540 15.335 -3.370 16.375 ;
        RECT -1.960 15.335 -1.790 16.375 ;
        RECT -0.380 15.335 -0.210 16.375 ;
        RECT 1.200 15.335 1.370 16.375 ;
        RECT 2.780 15.335 2.950 16.375 ;
        RECT 4.360 15.335 4.530 16.375 ;
        RECT 5.940 15.335 6.110 16.375 ;
        RECT 7.520 15.335 7.690 16.375 ;
        RECT 9.100 15.335 9.270 16.375 ;
        RECT 10.680 15.335 10.850 16.375 ;
        RECT -19.340 13.155 -19.170 14.195 ;
        RECT -17.760 13.155 -17.590 14.195 ;
        RECT -16.180 13.155 -16.010 14.195 ;
        RECT -14.600 13.155 -14.430 14.195 ;
        RECT -13.020 13.155 -12.850 14.195 ;
        RECT -11.440 13.155 -11.270 14.195 ;
        RECT -9.860 13.155 -9.690 14.195 ;
        RECT -8.280 13.155 -8.110 14.195 ;
        RECT -6.700 13.155 -6.530 14.195 ;
        RECT -5.120 13.155 -4.950 14.195 ;
        RECT -3.540 13.155 -3.370 14.195 ;
        RECT -1.960 13.155 -1.790 14.195 ;
        RECT -0.380 13.155 -0.210 14.195 ;
        RECT 1.200 13.155 1.370 14.195 ;
        RECT 2.780 13.155 2.950 14.195 ;
        RECT 4.360 13.155 4.530 14.195 ;
        RECT 5.940 13.155 6.110 14.195 ;
        RECT 7.520 13.155 7.690 14.195 ;
        RECT 9.100 13.155 9.270 14.195 ;
        RECT 10.680 13.155 10.850 14.195 ;
        RECT -19.340 10.975 -19.170 12.015 ;
        RECT -17.760 10.975 -17.590 12.015 ;
        RECT -16.180 10.975 -16.010 12.015 ;
        RECT -14.600 10.975 -14.430 12.015 ;
        RECT -13.020 10.975 -12.850 12.015 ;
        RECT -11.440 10.975 -11.270 12.015 ;
        RECT -9.860 10.975 -9.690 12.015 ;
        RECT -8.280 10.975 -8.110 12.015 ;
        RECT -6.700 10.975 -6.530 12.015 ;
        RECT -5.120 10.975 -4.950 12.015 ;
        RECT -3.540 10.975 -3.370 12.015 ;
        RECT -1.960 10.975 -1.790 12.015 ;
        RECT -0.380 10.975 -0.210 12.015 ;
        RECT 1.200 10.975 1.370 12.015 ;
        RECT 2.780 10.975 2.950 12.015 ;
        RECT 4.360 10.975 4.530 12.015 ;
        RECT 5.940 10.975 6.110 12.015 ;
        RECT 7.520 10.975 7.690 12.015 ;
        RECT 9.100 10.975 9.270 12.015 ;
        RECT 10.680 10.975 10.850 12.015 ;
        RECT -19.340 8.795 -19.170 9.835 ;
        RECT -17.760 8.795 -17.590 9.835 ;
        RECT -16.180 8.795 -16.010 9.835 ;
        RECT -14.600 8.795 -14.430 9.835 ;
        RECT -13.020 8.795 -12.850 9.835 ;
        RECT -11.440 8.795 -11.270 9.835 ;
        RECT -9.860 8.795 -9.690 9.835 ;
        RECT -8.280 8.795 -8.110 9.835 ;
        RECT -6.700 8.795 -6.530 9.835 ;
        RECT -5.120 8.795 -4.950 9.835 ;
        RECT -3.540 8.795 -3.370 9.835 ;
        RECT -1.960 8.795 -1.790 9.835 ;
        RECT -0.380 8.795 -0.210 9.835 ;
        RECT 1.200 8.795 1.370 9.835 ;
        RECT 2.780 8.795 2.950 9.835 ;
        RECT 4.360 8.795 4.530 9.835 ;
        RECT 5.940 8.795 6.110 9.835 ;
        RECT 7.520 8.795 7.690 9.835 ;
        RECT 9.100 8.795 9.270 9.835 ;
        RECT 10.680 8.795 10.850 9.835 ;
        RECT 12.140 7.890 13.655 19.445 ;
        RECT -22.305 5.885 13.655 7.890 ;
        RECT -22.305 4.950 -20.700 5.885 ;
        RECT -22.310 0.820 -20.700 4.950 ;
        RECT -17.475 4.770 13.655 5.885 ;
        RECT -17.475 2.270 -15.890 4.770 ;
        RECT -14.600 3.180 -14.430 4.220 ;
        RECT -13.140 2.270 -12.970 4.770 ;
        RECT -11.680 3.180 -11.510 4.220 ;
        RECT -10.220 2.270 -10.050 4.770 ;
        RECT -8.760 3.180 -8.590 4.220 ;
        RECT -7.300 2.270 -7.130 4.770 ;
        RECT -5.840 3.180 -5.670 4.220 ;
        RECT -4.380 2.270 -4.210 4.770 ;
        RECT -1.460 2.270 -1.290 4.770 ;
        RECT 1.460 2.270 1.630 4.770 ;
        RECT 2.920 3.180 3.090 4.220 ;
        RECT 4.380 2.270 4.550 4.770 ;
        RECT 5.050 3.180 5.220 4.220 ;
        RECT 6.510 2.270 8.050 4.770 ;
        RECT -17.475 1.815 8.050 2.270 ;
        RECT 11.870 0.940 13.655 4.770 ;
        RECT -22.310 -2.710 -21.480 0.820 ;
        RECT -22.305 -18.270 -21.480 -2.710 ;
        RECT 8.050 -16.950 10.210 -16.600 ;
        RECT 12.805 -18.270 13.655 0.940 ;
        RECT -22.305 -19.075 13.655 -18.270 ;
      LAYER met1 ;
        RECT -21.825 31.580 13.430 32.655 ;
        RECT -21.825 20.700 -21.170 31.580 ;
        RECT -19.370 29.650 -19.140 30.275 ;
        RECT -17.790 29.650 -17.560 30.275 ;
        RECT -16.210 29.650 -15.980 30.275 ;
        RECT -14.630 29.650 -14.400 30.275 ;
        RECT -13.050 29.650 -12.820 30.275 ;
        RECT -11.470 29.650 -11.240 30.275 ;
        RECT -9.890 29.650 -9.660 30.275 ;
        RECT -8.310 29.650 -8.080 30.275 ;
        RECT -6.730 29.650 -6.500 30.275 ;
        RECT -5.150 29.650 -4.920 30.275 ;
        RECT -3.570 29.650 -3.340 30.275 ;
        RECT -1.990 29.650 -1.760 30.275 ;
        RECT -0.410 29.650 -0.180 30.275 ;
        RECT 1.170 29.650 1.400 30.275 ;
        RECT 2.750 29.650 2.980 30.275 ;
        RECT 4.330 29.650 4.560 30.275 ;
        RECT 5.910 29.650 6.140 30.275 ;
        RECT 7.490 29.650 7.720 30.275 ;
        RECT 9.070 29.650 9.300 30.275 ;
        RECT 10.650 29.650 10.880 30.275 ;
        RECT -19.570 29.330 -18.930 29.650 ;
        RECT -17.990 29.330 -17.350 29.650 ;
        RECT -16.410 29.330 -15.770 29.650 ;
        RECT -14.830 29.330 -14.190 29.650 ;
        RECT -13.250 29.330 -12.610 29.650 ;
        RECT -11.670 29.330 -11.030 29.650 ;
        RECT -10.090 29.330 -9.450 29.650 ;
        RECT -8.510 29.330 -7.870 29.650 ;
        RECT -6.930 29.330 -6.290 29.650 ;
        RECT -5.350 29.330 -4.710 29.650 ;
        RECT -3.770 29.330 -3.130 29.650 ;
        RECT -2.190 29.330 -1.550 29.650 ;
        RECT -0.610 29.330 0.030 29.650 ;
        RECT 0.970 29.330 1.610 29.650 ;
        RECT 2.550 29.330 3.190 29.650 ;
        RECT 4.130 29.330 4.770 29.650 ;
        RECT 5.710 29.330 6.350 29.650 ;
        RECT 7.290 29.330 7.930 29.650 ;
        RECT 8.870 29.330 9.510 29.650 ;
        RECT 10.450 29.330 11.090 29.650 ;
        RECT -19.370 29.275 -19.140 29.330 ;
        RECT -17.790 29.275 -17.560 29.330 ;
        RECT -16.210 29.275 -15.980 29.330 ;
        RECT -14.630 29.275 -14.400 29.330 ;
        RECT -13.050 29.275 -12.820 29.330 ;
        RECT -11.470 29.275 -11.240 29.330 ;
        RECT -9.890 29.275 -9.660 29.330 ;
        RECT -8.310 29.275 -8.080 29.330 ;
        RECT -6.730 29.275 -6.500 29.330 ;
        RECT -5.150 29.275 -4.920 29.330 ;
        RECT -3.570 29.275 -3.340 29.330 ;
        RECT -1.990 29.275 -1.760 29.330 ;
        RECT -0.410 29.275 -0.180 29.330 ;
        RECT 1.170 29.275 1.400 29.330 ;
        RECT 2.750 29.275 2.980 29.330 ;
        RECT 4.330 29.275 4.560 29.330 ;
        RECT 5.910 29.275 6.140 29.330 ;
        RECT 7.490 29.275 7.720 29.330 ;
        RECT 9.070 29.275 9.300 29.330 ;
        RECT 10.650 29.275 10.880 29.330 ;
        RECT -19.370 27.450 -19.140 28.095 ;
        RECT -17.790 27.450 -17.560 28.095 ;
        RECT -16.210 27.450 -15.980 28.095 ;
        RECT -14.630 27.450 -14.400 28.095 ;
        RECT -13.050 27.450 -12.820 28.095 ;
        RECT -11.470 27.450 -11.240 28.095 ;
        RECT -9.890 27.450 -9.660 28.095 ;
        RECT -8.310 27.450 -8.080 28.095 ;
        RECT -6.730 27.450 -6.500 28.095 ;
        RECT -5.150 27.450 -4.920 28.095 ;
        RECT -3.570 27.450 -3.340 28.095 ;
        RECT -1.990 27.450 -1.760 28.095 ;
        RECT -0.410 27.450 -0.180 28.095 ;
        RECT 1.170 27.450 1.400 28.095 ;
        RECT 2.750 27.450 2.980 28.095 ;
        RECT 4.330 27.450 4.560 28.095 ;
        RECT 5.910 27.450 6.140 28.095 ;
        RECT 7.490 27.450 7.720 28.095 ;
        RECT 9.070 27.450 9.300 28.095 ;
        RECT 10.650 27.450 10.880 28.095 ;
        RECT -19.570 27.130 -18.930 27.450 ;
        RECT -17.990 27.130 -17.350 27.450 ;
        RECT -16.410 27.130 -15.770 27.450 ;
        RECT -14.830 27.130 -14.190 27.450 ;
        RECT -13.250 27.130 -12.610 27.450 ;
        RECT -11.670 27.130 -11.030 27.450 ;
        RECT -10.090 27.130 -9.450 27.450 ;
        RECT -8.510 27.130 -7.870 27.450 ;
        RECT -6.930 27.130 -6.290 27.450 ;
        RECT -5.350 27.130 -4.710 27.450 ;
        RECT -3.770 27.130 -3.130 27.450 ;
        RECT -2.190 27.130 -1.550 27.450 ;
        RECT -0.610 27.130 0.030 27.450 ;
        RECT 0.970 27.130 1.610 27.450 ;
        RECT 2.550 27.130 3.190 27.450 ;
        RECT 4.130 27.130 4.770 27.450 ;
        RECT 5.710 27.130 6.350 27.450 ;
        RECT 7.290 27.130 7.930 27.450 ;
        RECT 8.870 27.130 9.510 27.450 ;
        RECT 10.450 27.130 11.090 27.450 ;
        RECT -19.370 27.095 -19.140 27.130 ;
        RECT -17.790 27.095 -17.560 27.130 ;
        RECT -16.210 27.095 -15.980 27.130 ;
        RECT -14.630 27.095 -14.400 27.130 ;
        RECT -13.050 27.095 -12.820 27.130 ;
        RECT -11.470 27.095 -11.240 27.130 ;
        RECT -9.890 27.095 -9.660 27.130 ;
        RECT -8.310 27.095 -8.080 27.130 ;
        RECT -6.730 27.095 -6.500 27.130 ;
        RECT -5.150 27.095 -4.920 27.130 ;
        RECT -3.570 27.095 -3.340 27.130 ;
        RECT -1.990 27.095 -1.760 27.130 ;
        RECT -0.410 27.095 -0.180 27.130 ;
        RECT 1.170 27.095 1.400 27.130 ;
        RECT 2.750 27.095 2.980 27.130 ;
        RECT 4.330 27.095 4.560 27.130 ;
        RECT 5.910 27.095 6.140 27.130 ;
        RECT 7.490 27.095 7.720 27.130 ;
        RECT 9.070 27.095 9.300 27.130 ;
        RECT 10.650 27.095 10.880 27.130 ;
        RECT -19.370 25.250 -19.140 25.915 ;
        RECT -17.790 25.250 -17.560 25.915 ;
        RECT -16.210 25.250 -15.980 25.915 ;
        RECT -14.630 25.250 -14.400 25.915 ;
        RECT -13.050 25.250 -12.820 25.915 ;
        RECT -11.470 25.250 -11.240 25.915 ;
        RECT -9.890 25.250 -9.660 25.915 ;
        RECT -8.310 25.250 -8.080 25.915 ;
        RECT -6.730 25.250 -6.500 25.915 ;
        RECT -5.150 25.250 -4.920 25.915 ;
        RECT -3.570 25.250 -3.340 25.915 ;
        RECT -1.990 25.250 -1.760 25.915 ;
        RECT -0.410 25.250 -0.180 25.915 ;
        RECT 1.170 25.250 1.400 25.915 ;
        RECT 2.750 25.250 2.980 25.915 ;
        RECT 4.330 25.250 4.560 25.915 ;
        RECT 5.910 25.250 6.140 25.915 ;
        RECT 7.490 25.250 7.720 25.915 ;
        RECT 9.070 25.250 9.300 25.915 ;
        RECT 10.650 25.250 10.880 25.915 ;
        RECT -19.570 24.930 -18.930 25.250 ;
        RECT -17.990 24.930 -17.350 25.250 ;
        RECT -16.410 24.930 -15.770 25.250 ;
        RECT -14.830 24.930 -14.190 25.250 ;
        RECT -13.250 24.930 -12.610 25.250 ;
        RECT -11.670 24.930 -11.030 25.250 ;
        RECT -10.090 24.930 -9.450 25.250 ;
        RECT -8.510 24.930 -7.870 25.250 ;
        RECT -6.930 24.930 -6.290 25.250 ;
        RECT -5.350 24.930 -4.710 25.250 ;
        RECT -3.770 24.930 -3.130 25.250 ;
        RECT -2.190 24.930 -1.550 25.250 ;
        RECT -0.610 24.930 0.030 25.250 ;
        RECT 0.970 24.930 1.610 25.250 ;
        RECT 2.550 24.930 3.190 25.250 ;
        RECT 4.130 24.930 4.770 25.250 ;
        RECT 5.710 24.930 6.350 25.250 ;
        RECT 7.290 24.930 7.930 25.250 ;
        RECT 8.870 24.930 9.510 25.250 ;
        RECT 10.450 24.930 11.090 25.250 ;
        RECT -19.370 24.915 -19.140 24.930 ;
        RECT -17.790 24.915 -17.560 24.930 ;
        RECT -16.210 24.915 -15.980 24.930 ;
        RECT -14.630 24.915 -14.400 24.930 ;
        RECT -13.050 24.915 -12.820 24.930 ;
        RECT -11.470 24.915 -11.240 24.930 ;
        RECT -9.890 24.915 -9.660 24.930 ;
        RECT -8.310 24.915 -8.080 24.930 ;
        RECT -6.730 24.915 -6.500 24.930 ;
        RECT -5.150 24.915 -4.920 24.930 ;
        RECT -3.570 24.915 -3.340 24.930 ;
        RECT -1.990 24.915 -1.760 24.930 ;
        RECT -0.410 24.915 -0.180 24.930 ;
        RECT 1.170 24.915 1.400 24.930 ;
        RECT 2.750 24.915 2.980 24.930 ;
        RECT 4.330 24.915 4.560 24.930 ;
        RECT 5.910 24.915 6.140 24.930 ;
        RECT 7.490 24.915 7.720 24.930 ;
        RECT 9.070 24.915 9.300 24.930 ;
        RECT 10.650 24.915 10.880 24.930 ;
        RECT -19.370 23.075 -19.140 23.735 ;
        RECT -17.790 23.075 -17.560 23.735 ;
        RECT -16.210 23.075 -15.980 23.735 ;
        RECT -14.630 23.075 -14.400 23.735 ;
        RECT -13.050 23.075 -12.820 23.735 ;
        RECT -11.470 23.075 -11.240 23.735 ;
        RECT -9.890 23.075 -9.660 23.735 ;
        RECT -8.310 23.075 -8.080 23.735 ;
        RECT -6.730 23.075 -6.500 23.735 ;
        RECT -5.150 23.075 -4.920 23.735 ;
        RECT -3.570 23.075 -3.340 23.735 ;
        RECT -1.990 23.075 -1.760 23.735 ;
        RECT -0.410 23.075 -0.180 23.735 ;
        RECT 1.170 23.075 1.400 23.735 ;
        RECT 2.750 23.075 2.980 23.735 ;
        RECT 4.330 23.075 4.560 23.735 ;
        RECT 5.910 23.075 6.140 23.735 ;
        RECT 7.490 23.075 7.720 23.735 ;
        RECT 9.070 23.075 9.300 23.735 ;
        RECT 10.650 23.075 10.880 23.735 ;
        RECT -19.570 22.755 -18.930 23.075 ;
        RECT -17.990 22.755 -17.350 23.075 ;
        RECT -16.410 22.755 -15.770 23.075 ;
        RECT -14.830 22.755 -14.190 23.075 ;
        RECT -13.250 22.755 -12.610 23.075 ;
        RECT -11.670 22.755 -11.030 23.075 ;
        RECT -10.090 22.755 -9.450 23.075 ;
        RECT -8.510 22.755 -7.870 23.075 ;
        RECT -6.930 22.755 -6.290 23.075 ;
        RECT -5.350 22.755 -4.710 23.075 ;
        RECT -3.770 22.755 -3.130 23.075 ;
        RECT -2.190 22.755 -1.550 23.075 ;
        RECT -0.610 22.755 0.030 23.075 ;
        RECT 0.970 22.755 1.610 23.075 ;
        RECT 2.550 22.755 3.190 23.075 ;
        RECT 4.130 22.755 4.770 23.075 ;
        RECT 5.710 22.755 6.350 23.075 ;
        RECT 7.290 22.755 7.930 23.075 ;
        RECT 8.870 22.755 9.510 23.075 ;
        RECT 10.450 22.755 11.090 23.075 ;
        RECT -19.370 22.735 -19.140 22.755 ;
        RECT -17.790 22.735 -17.560 22.755 ;
        RECT -16.210 22.735 -15.980 22.755 ;
        RECT -14.630 22.735 -14.400 22.755 ;
        RECT -13.050 22.735 -12.820 22.755 ;
        RECT -11.470 22.735 -11.240 22.755 ;
        RECT -9.890 22.735 -9.660 22.755 ;
        RECT -8.310 22.735 -8.080 22.755 ;
        RECT -6.730 22.735 -6.500 22.755 ;
        RECT -5.150 22.735 -4.920 22.755 ;
        RECT -3.570 22.735 -3.340 22.755 ;
        RECT -1.990 22.735 -1.760 22.755 ;
        RECT -0.410 22.735 -0.180 22.755 ;
        RECT 1.170 22.735 1.400 22.755 ;
        RECT 2.750 22.735 2.980 22.755 ;
        RECT 4.330 22.735 4.560 22.755 ;
        RECT 5.910 22.735 6.140 22.755 ;
        RECT 7.490 22.735 7.720 22.755 ;
        RECT 9.070 22.735 9.300 22.755 ;
        RECT 10.650 22.735 10.880 22.755 ;
        RECT -19.370 20.950 -19.140 21.555 ;
        RECT -17.790 20.950 -17.560 21.555 ;
        RECT -16.210 20.950 -15.980 21.555 ;
        RECT -14.630 20.950 -14.400 21.555 ;
        RECT -13.050 20.950 -12.820 21.555 ;
        RECT -11.470 20.950 -11.240 21.555 ;
        RECT -9.890 20.950 -9.660 21.555 ;
        RECT -8.310 20.950 -8.080 21.555 ;
        RECT -6.730 20.950 -6.500 21.555 ;
        RECT -5.150 20.950 -4.920 21.555 ;
        RECT -3.570 20.950 -3.340 21.555 ;
        RECT -1.990 20.950 -1.760 21.555 ;
        RECT -0.410 20.950 -0.180 21.555 ;
        RECT 1.170 20.950 1.400 21.555 ;
        RECT 2.750 20.950 2.980 21.555 ;
        RECT 4.330 20.950 4.560 21.555 ;
        RECT 5.910 20.950 6.140 21.555 ;
        RECT 7.490 20.950 7.720 21.555 ;
        RECT 9.070 20.950 9.300 21.555 ;
        RECT 10.650 20.950 10.880 21.555 ;
        RECT -19.570 20.630 -18.930 20.950 ;
        RECT -17.990 20.630 -17.350 20.950 ;
        RECT -16.410 20.630 -15.770 20.950 ;
        RECT -14.830 20.630 -14.190 20.950 ;
        RECT -13.250 20.630 -12.610 20.950 ;
        RECT -11.670 20.630 -11.030 20.950 ;
        RECT -10.090 20.630 -9.450 20.950 ;
        RECT -8.510 20.630 -7.870 20.950 ;
        RECT -6.930 20.630 -6.290 20.950 ;
        RECT -5.350 20.630 -4.710 20.950 ;
        RECT -3.770 20.630 -3.130 20.950 ;
        RECT -2.190 20.630 -1.550 20.950 ;
        RECT -0.610 20.630 0.030 20.950 ;
        RECT 0.970 20.630 1.610 20.950 ;
        RECT 2.550 20.630 3.190 20.950 ;
        RECT 4.130 20.630 4.770 20.950 ;
        RECT 5.710 20.630 6.350 20.950 ;
        RECT 7.290 20.630 7.930 20.950 ;
        RECT 8.870 20.630 9.510 20.950 ;
        RECT 10.450 20.630 11.090 20.950 ;
        RECT -19.370 20.555 -19.140 20.630 ;
        RECT -17.790 20.555 -17.560 20.630 ;
        RECT -16.210 20.555 -15.980 20.630 ;
        RECT -14.630 20.555 -14.400 20.630 ;
        RECT -13.050 20.555 -12.820 20.630 ;
        RECT -11.470 20.555 -11.240 20.630 ;
        RECT -9.890 20.555 -9.660 20.630 ;
        RECT -8.310 20.555 -8.080 20.630 ;
        RECT -6.730 20.555 -6.500 20.630 ;
        RECT -5.150 20.555 -4.920 20.630 ;
        RECT -3.570 20.555 -3.340 20.630 ;
        RECT -1.990 20.555 -1.760 20.630 ;
        RECT -0.410 20.555 -0.180 20.630 ;
        RECT 1.170 20.555 1.400 20.630 ;
        RECT 2.750 20.555 2.980 20.630 ;
        RECT 4.330 20.555 4.560 20.630 ;
        RECT 5.910 20.555 6.140 20.630 ;
        RECT 7.490 20.555 7.720 20.630 ;
        RECT 9.070 20.555 9.300 20.630 ;
        RECT 10.650 20.555 10.880 20.630 ;
        RECT -20.850 19.405 12.425 19.705 ;
        RECT -19.370 17.850 -19.140 18.535 ;
        RECT -17.790 17.850 -17.560 18.535 ;
        RECT -16.210 17.850 -15.980 18.535 ;
        RECT -14.630 17.850 -14.400 18.535 ;
        RECT -13.050 17.850 -12.820 18.535 ;
        RECT -11.470 17.850 -11.240 18.535 ;
        RECT -9.890 17.850 -9.660 18.535 ;
        RECT -8.310 17.850 -8.080 18.535 ;
        RECT -6.730 17.850 -6.500 18.535 ;
        RECT -5.150 17.850 -4.920 18.535 ;
        RECT -3.570 17.850 -3.340 18.535 ;
        RECT -1.990 17.850 -1.760 18.535 ;
        RECT -0.410 17.850 -0.180 18.535 ;
        RECT 1.170 17.850 1.400 18.535 ;
        RECT 2.750 17.850 2.980 18.535 ;
        RECT 4.330 17.850 4.560 18.535 ;
        RECT 5.910 17.850 6.140 18.535 ;
        RECT 7.490 17.850 7.720 18.535 ;
        RECT 9.070 17.850 9.300 18.535 ;
        RECT 10.650 17.850 10.880 18.535 ;
        RECT -19.570 17.530 -18.930 17.850 ;
        RECT -17.990 17.530 -17.350 17.850 ;
        RECT -16.410 17.530 -15.770 17.850 ;
        RECT -14.830 17.530 -14.190 17.850 ;
        RECT -13.250 17.530 -12.610 17.850 ;
        RECT -11.670 17.530 -11.030 17.850 ;
        RECT -10.090 17.530 -9.450 17.850 ;
        RECT -8.510 17.530 -7.870 17.850 ;
        RECT -6.930 17.530 -6.290 17.850 ;
        RECT -5.350 17.530 -4.710 17.850 ;
        RECT -3.770 17.530 -3.130 17.850 ;
        RECT -2.190 17.530 -1.550 17.850 ;
        RECT -0.610 17.530 0.030 17.850 ;
        RECT 0.970 17.530 1.610 17.850 ;
        RECT 2.550 17.530 3.190 17.850 ;
        RECT 4.130 17.530 4.770 17.850 ;
        RECT 5.710 17.530 6.350 17.850 ;
        RECT 7.290 17.530 7.930 17.850 ;
        RECT 8.870 17.530 9.510 17.850 ;
        RECT 10.450 17.530 11.090 17.850 ;
        RECT -19.370 15.675 -19.140 16.355 ;
        RECT -17.790 15.675 -17.560 16.355 ;
        RECT -16.210 15.675 -15.980 16.355 ;
        RECT -14.630 15.675 -14.400 16.355 ;
        RECT -13.050 15.675 -12.820 16.355 ;
        RECT -11.470 15.675 -11.240 16.355 ;
        RECT -9.890 15.675 -9.660 16.355 ;
        RECT -8.310 15.675 -8.080 16.355 ;
        RECT -6.730 15.675 -6.500 16.355 ;
        RECT -5.150 15.675 -4.920 16.355 ;
        RECT -3.570 15.675 -3.340 16.355 ;
        RECT -1.990 15.675 -1.760 16.355 ;
        RECT -0.410 15.675 -0.180 16.355 ;
        RECT 1.170 15.675 1.400 16.355 ;
        RECT 2.750 15.675 2.980 16.355 ;
        RECT 4.330 15.675 4.560 16.355 ;
        RECT 5.910 15.675 6.140 16.355 ;
        RECT 7.490 15.675 7.720 16.355 ;
        RECT 9.070 15.675 9.300 16.355 ;
        RECT 10.650 15.675 10.880 16.355 ;
        RECT -19.570 15.355 -18.930 15.675 ;
        RECT -17.990 15.355 -17.350 15.675 ;
        RECT -16.410 15.355 -15.770 15.675 ;
        RECT -14.830 15.355 -14.190 15.675 ;
        RECT -13.250 15.355 -12.610 15.675 ;
        RECT -11.670 15.355 -11.030 15.675 ;
        RECT -10.090 15.355 -9.450 15.675 ;
        RECT -8.510 15.355 -7.870 15.675 ;
        RECT -6.930 15.355 -6.290 15.675 ;
        RECT -5.350 15.355 -4.710 15.675 ;
        RECT -3.770 15.355 -3.130 15.675 ;
        RECT -2.190 15.355 -1.550 15.675 ;
        RECT -0.610 15.355 0.030 15.675 ;
        RECT 0.970 15.355 1.610 15.675 ;
        RECT 2.550 15.355 3.190 15.675 ;
        RECT 4.130 15.355 4.770 15.675 ;
        RECT 5.710 15.355 6.350 15.675 ;
        RECT 7.290 15.355 7.930 15.675 ;
        RECT 8.870 15.355 9.510 15.675 ;
        RECT 10.450 15.355 11.090 15.675 ;
        RECT -19.370 13.500 -19.140 14.175 ;
        RECT -17.790 13.500 -17.560 14.175 ;
        RECT -16.210 13.500 -15.980 14.175 ;
        RECT -14.630 13.500 -14.400 14.175 ;
        RECT -13.050 13.500 -12.820 14.175 ;
        RECT -11.470 13.500 -11.240 14.175 ;
        RECT -9.890 13.500 -9.660 14.175 ;
        RECT -8.310 13.500 -8.080 14.175 ;
        RECT -6.730 13.500 -6.500 14.175 ;
        RECT -5.150 13.500 -4.920 14.175 ;
        RECT -3.570 13.500 -3.340 14.175 ;
        RECT -1.990 13.500 -1.760 14.175 ;
        RECT -0.410 13.500 -0.180 14.175 ;
        RECT 1.170 13.500 1.400 14.175 ;
        RECT 2.750 13.500 2.980 14.175 ;
        RECT 4.330 13.500 4.560 14.175 ;
        RECT 5.910 13.500 6.140 14.175 ;
        RECT 7.490 13.500 7.720 14.175 ;
        RECT 9.070 13.500 9.300 14.175 ;
        RECT 10.650 13.500 10.880 14.175 ;
        RECT -19.570 13.180 -18.930 13.500 ;
        RECT -17.990 13.180 -17.350 13.500 ;
        RECT -16.410 13.180 -15.770 13.500 ;
        RECT -14.830 13.180 -14.190 13.500 ;
        RECT -13.250 13.180 -12.610 13.500 ;
        RECT -11.670 13.180 -11.030 13.500 ;
        RECT -10.090 13.180 -9.450 13.500 ;
        RECT -8.510 13.180 -7.870 13.500 ;
        RECT -6.930 13.180 -6.290 13.500 ;
        RECT -5.350 13.180 -4.710 13.500 ;
        RECT -3.770 13.180 -3.130 13.500 ;
        RECT -2.190 13.180 -1.550 13.500 ;
        RECT -0.610 13.180 0.030 13.500 ;
        RECT 0.970 13.180 1.610 13.500 ;
        RECT 2.550 13.180 3.190 13.500 ;
        RECT 4.130 13.180 4.770 13.500 ;
        RECT 5.710 13.180 6.350 13.500 ;
        RECT 7.290 13.180 7.930 13.500 ;
        RECT 8.870 13.180 9.510 13.500 ;
        RECT 10.450 13.180 11.090 13.500 ;
        RECT -19.370 13.175 -19.140 13.180 ;
        RECT -17.790 13.175 -17.560 13.180 ;
        RECT -16.210 13.175 -15.980 13.180 ;
        RECT -14.630 13.175 -14.400 13.180 ;
        RECT -13.050 13.175 -12.820 13.180 ;
        RECT -11.470 13.175 -11.240 13.180 ;
        RECT -9.890 13.175 -9.660 13.180 ;
        RECT -8.310 13.175 -8.080 13.180 ;
        RECT -6.730 13.175 -6.500 13.180 ;
        RECT -5.150 13.175 -4.920 13.180 ;
        RECT -3.570 13.175 -3.340 13.180 ;
        RECT -1.990 13.175 -1.760 13.180 ;
        RECT -0.410 13.175 -0.180 13.180 ;
        RECT 1.170 13.175 1.400 13.180 ;
        RECT 2.750 13.175 2.980 13.180 ;
        RECT 4.330 13.175 4.560 13.180 ;
        RECT 5.910 13.175 6.140 13.180 ;
        RECT 7.490 13.175 7.720 13.180 ;
        RECT 9.070 13.175 9.300 13.180 ;
        RECT 10.650 13.175 10.880 13.180 ;
        RECT -19.370 11.325 -19.140 11.995 ;
        RECT -17.790 11.325 -17.560 11.995 ;
        RECT -16.210 11.325 -15.980 11.995 ;
        RECT -14.630 11.325 -14.400 11.995 ;
        RECT -13.050 11.325 -12.820 11.995 ;
        RECT -11.470 11.325 -11.240 11.995 ;
        RECT -9.890 11.325 -9.660 11.995 ;
        RECT -8.310 11.325 -8.080 11.995 ;
        RECT -6.730 11.325 -6.500 11.995 ;
        RECT -5.150 11.325 -4.920 11.995 ;
        RECT -3.570 11.325 -3.340 11.995 ;
        RECT -1.990 11.325 -1.760 11.995 ;
        RECT -0.410 11.325 -0.180 11.995 ;
        RECT 1.170 11.325 1.400 11.995 ;
        RECT 2.750 11.325 2.980 11.995 ;
        RECT 4.330 11.325 4.560 11.995 ;
        RECT 5.910 11.325 6.140 11.995 ;
        RECT 7.490 11.325 7.720 11.995 ;
        RECT 9.070 11.325 9.300 11.995 ;
        RECT 10.650 11.325 10.880 11.995 ;
        RECT -19.570 11.005 -18.930 11.325 ;
        RECT -17.990 11.005 -17.350 11.325 ;
        RECT -16.410 11.005 -15.770 11.325 ;
        RECT -14.830 11.005 -14.190 11.325 ;
        RECT -13.250 11.005 -12.610 11.325 ;
        RECT -11.670 11.005 -11.030 11.325 ;
        RECT -10.090 11.005 -9.450 11.325 ;
        RECT -8.510 11.005 -7.870 11.325 ;
        RECT -6.930 11.005 -6.290 11.325 ;
        RECT -5.350 11.005 -4.710 11.325 ;
        RECT -3.770 11.005 -3.130 11.325 ;
        RECT -2.190 11.005 -1.550 11.325 ;
        RECT -0.610 11.005 0.030 11.325 ;
        RECT 0.970 11.005 1.610 11.325 ;
        RECT 2.550 11.005 3.190 11.325 ;
        RECT 4.130 11.005 4.770 11.325 ;
        RECT 5.710 11.005 6.350 11.325 ;
        RECT 7.290 11.005 7.930 11.325 ;
        RECT 8.870 11.005 9.510 11.325 ;
        RECT 10.450 11.005 11.090 11.325 ;
        RECT -19.370 10.995 -19.140 11.005 ;
        RECT -17.790 10.995 -17.560 11.005 ;
        RECT -16.210 10.995 -15.980 11.005 ;
        RECT -14.630 10.995 -14.400 11.005 ;
        RECT -13.050 10.995 -12.820 11.005 ;
        RECT -11.470 10.995 -11.240 11.005 ;
        RECT -9.890 10.995 -9.660 11.005 ;
        RECT -8.310 10.995 -8.080 11.005 ;
        RECT -6.730 10.995 -6.500 11.005 ;
        RECT -5.150 10.995 -4.920 11.005 ;
        RECT -3.570 10.995 -3.340 11.005 ;
        RECT -1.990 10.995 -1.760 11.005 ;
        RECT -0.410 10.995 -0.180 11.005 ;
        RECT 1.170 10.995 1.400 11.005 ;
        RECT 2.750 10.995 2.980 11.005 ;
        RECT 4.330 10.995 4.560 11.005 ;
        RECT 5.910 10.995 6.140 11.005 ;
        RECT 7.490 10.995 7.720 11.005 ;
        RECT 9.070 10.995 9.300 11.005 ;
        RECT 10.650 10.995 10.880 11.005 ;
        RECT -19.370 9.150 -19.140 9.815 ;
        RECT -17.790 9.150 -17.560 9.815 ;
        RECT -16.210 9.150 -15.980 9.815 ;
        RECT -14.630 9.150 -14.400 9.815 ;
        RECT -13.050 9.150 -12.820 9.815 ;
        RECT -11.470 9.150 -11.240 9.815 ;
        RECT -9.890 9.150 -9.660 9.815 ;
        RECT -8.310 9.150 -8.080 9.815 ;
        RECT -6.730 9.150 -6.500 9.815 ;
        RECT -5.150 9.150 -4.920 9.815 ;
        RECT -3.570 9.150 -3.340 9.815 ;
        RECT -1.990 9.150 -1.760 9.815 ;
        RECT -0.410 9.150 -0.180 9.815 ;
        RECT 1.170 9.150 1.400 9.815 ;
        RECT 2.750 9.150 2.980 9.815 ;
        RECT 4.330 9.150 4.560 9.815 ;
        RECT 5.910 9.150 6.140 9.815 ;
        RECT 7.490 9.150 7.720 9.815 ;
        RECT 9.070 9.150 9.300 9.815 ;
        RECT 10.650 9.150 10.880 9.815 ;
        RECT -19.570 8.830 -18.930 9.150 ;
        RECT -17.990 8.830 -17.350 9.150 ;
        RECT -16.410 8.830 -15.770 9.150 ;
        RECT -14.830 8.830 -14.190 9.150 ;
        RECT -13.250 8.830 -12.610 9.150 ;
        RECT -11.670 8.830 -11.030 9.150 ;
        RECT -10.090 8.830 -9.450 9.150 ;
        RECT -8.510 8.830 -7.870 9.150 ;
        RECT -6.930 8.830 -6.290 9.150 ;
        RECT -5.350 8.830 -4.710 9.150 ;
        RECT -3.770 8.830 -3.130 9.150 ;
        RECT -2.190 8.830 -1.550 9.150 ;
        RECT -0.610 8.830 0.030 9.150 ;
        RECT 0.970 8.830 1.610 9.150 ;
        RECT 2.550 8.830 3.190 9.150 ;
        RECT 4.130 8.830 4.770 9.150 ;
        RECT 5.710 8.830 6.350 9.150 ;
        RECT 7.290 8.830 7.930 9.150 ;
        RECT 8.870 8.830 9.510 9.150 ;
        RECT 10.450 8.830 11.090 9.150 ;
        RECT -19.370 8.815 -19.140 8.830 ;
        RECT -17.790 8.815 -17.560 8.830 ;
        RECT -16.210 8.815 -15.980 8.830 ;
        RECT -14.630 8.815 -14.400 8.830 ;
        RECT -13.050 8.815 -12.820 8.830 ;
        RECT -11.470 8.815 -11.240 8.830 ;
        RECT -9.890 8.815 -9.660 8.830 ;
        RECT -8.310 8.815 -8.080 8.830 ;
        RECT -6.730 8.815 -6.500 8.830 ;
        RECT -5.150 8.815 -4.920 8.830 ;
        RECT -3.570 8.815 -3.340 8.830 ;
        RECT -1.990 8.815 -1.760 8.830 ;
        RECT -0.410 8.815 -0.180 8.830 ;
        RECT 1.170 8.815 1.400 8.830 ;
        RECT 2.750 8.815 2.980 8.830 ;
        RECT 4.330 8.815 4.560 8.830 ;
        RECT 5.910 8.815 6.140 8.830 ;
        RECT 7.490 8.815 7.720 8.830 ;
        RECT 9.070 8.815 9.300 8.830 ;
        RECT 10.650 8.815 10.880 8.830 ;
        RECT -21.810 5.530 -20.700 7.005 ;
        RECT -20.385 5.885 -19.065 7.225 ;
        RECT -17.220 5.905 7.765 7.245 ;
        RECT -17.220 2.990 -16.230 5.905 ;
        RECT -14.735 5.885 -5.495 5.905 ;
        RECT 2.235 5.885 3.745 5.905 ;
        RECT -14.735 3.200 -14.270 5.885 ;
        RECT -11.780 3.190 -11.315 5.885 ;
        RECT -8.895 3.180 -8.430 5.885 ;
        RECT -5.960 3.190 -5.495 5.885 ;
        RECT 2.695 3.200 3.335 5.885 ;
        RECT 5.020 4.140 5.250 4.200 ;
        RECT 4.930 3.260 5.365 4.140 ;
        RECT 5.020 3.200 5.250 3.260 ;
        RECT 6.865 2.305 7.765 5.905 ;
        RECT 10.555 5.455 13.415 7.225 ;
        RECT 10.555 -1.065 11.815 5.455 ;
        RECT 10.555 -1.415 13.495 -1.065 ;
        RECT -22.170 -10.275 -21.480 -3.035 ;
        RECT 13.145 -12.345 13.495 -1.415 ;
        RECT -22.170 -18.270 -21.480 -12.740 ;
        RECT 7.990 -17.330 11.140 -16.195 ;
        RECT 12.805 -18.270 13.495 -12.345 ;
        RECT -22.170 -18.960 13.495 -18.270 ;
      LAYER met2 ;
        RECT -21.810 31.565 13.425 32.675 ;
        RECT -21.810 29.655 -20.700 31.565 ;
        RECT -21.810 29.650 -20.405 29.655 ;
        RECT -21.810 28.960 11.995 29.650 ;
        RECT -21.810 27.450 -20.700 28.960 ;
        RECT -20.405 28.955 11.995 28.960 ;
        RECT -21.810 26.755 11.995 27.450 ;
        RECT -21.810 25.250 -20.700 26.755 ;
        RECT -21.810 24.555 11.995 25.250 ;
        RECT -21.810 23.075 -20.700 24.555 ;
        RECT -21.810 22.380 11.995 23.075 ;
        RECT -21.810 20.950 -20.700 22.380 ;
        RECT -21.810 20.255 11.995 20.950 ;
        RECT -21.810 19.705 -20.700 20.255 ;
        RECT -21.810 19.405 11.880 19.705 ;
        RECT -21.810 17.850 -20.700 19.405 ;
        RECT -21.810 17.155 11.995 17.850 ;
        RECT -21.810 15.675 -20.700 17.155 ;
        RECT -21.810 14.980 11.995 15.675 ;
        RECT -21.810 13.500 -20.700 14.980 ;
        RECT -21.810 12.805 11.995 13.500 ;
        RECT -21.810 11.325 -20.700 12.805 ;
        RECT -21.810 10.630 11.995 11.325 ;
        RECT -21.810 9.150 -20.700 10.630 ;
        RECT -21.810 8.455 11.995 9.150 ;
        RECT -27.390 7.010 -25.700 7.240 ;
        RECT -21.810 7.225 -20.700 8.455 ;
        RECT -21.810 7.010 11.815 7.225 ;
        RECT -27.390 6.000 11.815 7.010 ;
        RECT -27.390 5.650 -25.700 6.000 ;
        RECT -21.810 5.885 11.815 6.000 ;
        RECT -21.810 5.530 -20.700 5.885 ;
        RECT 4.885 3.260 5.410 5.885 ;
        RECT 7.865 -17.455 13.525 -16.100 ;
      LAYER met3 ;
        RECT -27.300 5.785 -25.850 7.135 ;
      LAYER met4 ;
        RECT -27.390 33.300 16.870 34.950 ;
        RECT -27.255 5.805 -25.895 7.115 ;
        RECT -27.390 -21.200 16.870 -19.550 ;
      LAYER met5 ;
        RECT -27.390 33.170 -25.710 34.950 ;
        RECT 15.160 33.310 16.860 34.950 ;
        RECT -27.390 -20.550 -25.700 33.170 ;
        RECT -27.390 -21.200 -25.710 -20.550 ;
        RECT 15.160 -21.200 16.840 33.310 ;
    END
  END vdd
  PIN out
    ANTENNADIFFAREA 79.169998 ;
    PORT
      LAYER li1 ;
        RECT -20.130 29.255 -19.960 30.295 ;
        RECT -18.550 29.255 -18.380 30.295 ;
        RECT -16.970 29.255 -16.800 30.295 ;
        RECT -15.390 29.255 -15.220 30.295 ;
        RECT -13.810 29.255 -13.640 30.295 ;
        RECT -12.230 29.255 -12.060 30.295 ;
        RECT -10.650 29.255 -10.480 30.295 ;
        RECT -9.070 29.255 -8.900 30.295 ;
        RECT -7.490 29.255 -7.320 30.295 ;
        RECT -5.910 29.255 -5.740 30.295 ;
        RECT -4.330 29.255 -4.160 30.295 ;
        RECT -2.750 29.255 -2.580 30.295 ;
        RECT -1.170 29.255 -1.000 30.295 ;
        RECT 0.410 29.255 0.580 30.295 ;
        RECT 1.990 29.255 2.160 30.295 ;
        RECT 3.570 29.255 3.740 30.295 ;
        RECT 5.150 29.255 5.320 30.295 ;
        RECT 6.730 29.255 6.900 30.295 ;
        RECT 8.310 29.255 8.480 30.295 ;
        RECT 9.890 29.255 10.060 30.295 ;
        RECT 11.470 29.255 11.640 30.295 ;
        RECT -20.130 27.075 -19.960 28.115 ;
        RECT -18.550 27.075 -18.380 28.115 ;
        RECT -16.970 27.075 -16.800 28.115 ;
        RECT -15.390 27.075 -15.220 28.115 ;
        RECT -13.810 27.075 -13.640 28.115 ;
        RECT -12.230 27.075 -12.060 28.115 ;
        RECT -10.650 27.075 -10.480 28.115 ;
        RECT -9.070 27.075 -8.900 28.115 ;
        RECT -7.490 27.075 -7.320 28.115 ;
        RECT -5.910 27.075 -5.740 28.115 ;
        RECT -4.330 27.075 -4.160 28.115 ;
        RECT -2.750 27.075 -2.580 28.115 ;
        RECT -1.170 27.075 -1.000 28.115 ;
        RECT 0.410 27.075 0.580 28.115 ;
        RECT 1.990 27.075 2.160 28.115 ;
        RECT 3.570 27.075 3.740 28.115 ;
        RECT 5.150 27.075 5.320 28.115 ;
        RECT 6.730 27.075 6.900 28.115 ;
        RECT 8.310 27.075 8.480 28.115 ;
        RECT 9.890 27.075 10.060 28.115 ;
        RECT 11.470 27.075 11.640 28.115 ;
        RECT -20.130 24.895 -19.960 25.935 ;
        RECT -18.550 24.895 -18.380 25.935 ;
        RECT -16.970 24.895 -16.800 25.935 ;
        RECT -15.390 24.895 -15.220 25.935 ;
        RECT -13.810 24.895 -13.640 25.935 ;
        RECT -12.230 24.895 -12.060 25.935 ;
        RECT -10.650 24.895 -10.480 25.935 ;
        RECT -9.070 24.895 -8.900 25.935 ;
        RECT -7.490 24.895 -7.320 25.935 ;
        RECT -5.910 24.895 -5.740 25.935 ;
        RECT -4.330 24.895 -4.160 25.935 ;
        RECT -2.750 24.895 -2.580 25.935 ;
        RECT -1.170 24.895 -1.000 25.935 ;
        RECT 0.410 24.895 0.580 25.935 ;
        RECT 1.990 24.895 2.160 25.935 ;
        RECT 3.570 24.895 3.740 25.935 ;
        RECT 5.150 24.895 5.320 25.935 ;
        RECT 6.730 24.895 6.900 25.935 ;
        RECT 8.310 24.895 8.480 25.935 ;
        RECT 9.890 24.895 10.060 25.935 ;
        RECT 11.470 24.895 11.640 25.935 ;
        RECT -20.130 22.715 -19.960 23.755 ;
        RECT -18.550 22.715 -18.380 23.755 ;
        RECT -16.970 22.715 -16.800 23.755 ;
        RECT -15.390 22.715 -15.220 23.755 ;
        RECT -13.810 22.715 -13.640 23.755 ;
        RECT -12.230 22.715 -12.060 23.755 ;
        RECT -10.650 22.715 -10.480 23.755 ;
        RECT -9.070 22.715 -8.900 23.755 ;
        RECT -7.490 22.715 -7.320 23.755 ;
        RECT -5.910 22.715 -5.740 23.755 ;
        RECT -4.330 22.715 -4.160 23.755 ;
        RECT -2.750 22.715 -2.580 23.755 ;
        RECT -1.170 22.715 -1.000 23.755 ;
        RECT 0.410 22.715 0.580 23.755 ;
        RECT 1.990 22.715 2.160 23.755 ;
        RECT 3.570 22.715 3.740 23.755 ;
        RECT 5.150 22.715 5.320 23.755 ;
        RECT 6.730 22.715 6.900 23.755 ;
        RECT 8.310 22.715 8.480 23.755 ;
        RECT 9.890 22.715 10.060 23.755 ;
        RECT 11.470 22.715 11.640 23.755 ;
        RECT -20.130 20.535 -19.960 21.575 ;
        RECT -18.550 20.535 -18.380 21.575 ;
        RECT -16.970 20.535 -16.800 21.575 ;
        RECT -15.390 20.535 -15.220 21.575 ;
        RECT -13.810 20.535 -13.640 21.575 ;
        RECT -12.230 20.535 -12.060 21.575 ;
        RECT -10.650 20.535 -10.480 21.575 ;
        RECT -9.070 20.535 -8.900 21.575 ;
        RECT -7.490 20.535 -7.320 21.575 ;
        RECT -5.910 20.535 -5.740 21.575 ;
        RECT -4.330 20.535 -4.160 21.575 ;
        RECT -2.750 20.535 -2.580 21.575 ;
        RECT -1.170 20.535 -1.000 21.575 ;
        RECT 0.410 20.535 0.580 21.575 ;
        RECT 1.990 20.535 2.160 21.575 ;
        RECT 3.570 20.535 3.740 21.575 ;
        RECT 5.150 20.535 5.320 21.575 ;
        RECT 6.730 20.535 6.900 21.575 ;
        RECT 8.310 20.535 8.480 21.575 ;
        RECT 9.890 20.535 10.060 21.575 ;
        RECT 11.470 20.535 11.640 21.575 ;
        RECT -20.130 17.515 -19.960 18.555 ;
        RECT -18.550 17.515 -18.380 18.555 ;
        RECT -16.970 17.515 -16.800 18.555 ;
        RECT -15.390 17.515 -15.220 18.555 ;
        RECT -13.810 17.515 -13.640 18.555 ;
        RECT -12.230 17.515 -12.060 18.555 ;
        RECT -10.650 17.515 -10.480 18.555 ;
        RECT -9.070 17.515 -8.900 18.555 ;
        RECT -7.490 17.515 -7.320 18.555 ;
        RECT -5.910 17.515 -5.740 18.555 ;
        RECT -4.330 17.515 -4.160 18.555 ;
        RECT -2.750 17.515 -2.580 18.555 ;
        RECT -1.170 17.515 -1.000 18.555 ;
        RECT 0.410 17.515 0.580 18.555 ;
        RECT 1.990 17.515 2.160 18.555 ;
        RECT 3.570 17.515 3.740 18.555 ;
        RECT 5.150 17.515 5.320 18.555 ;
        RECT 6.730 17.515 6.900 18.555 ;
        RECT 8.310 17.515 8.480 18.555 ;
        RECT 9.890 17.515 10.060 18.555 ;
        RECT 11.470 17.515 11.640 18.555 ;
        RECT -20.130 15.335 -19.960 16.375 ;
        RECT -18.550 15.335 -18.380 16.375 ;
        RECT -16.970 15.335 -16.800 16.375 ;
        RECT -15.390 15.335 -15.220 16.375 ;
        RECT -13.810 15.335 -13.640 16.375 ;
        RECT -12.230 15.335 -12.060 16.375 ;
        RECT -10.650 15.335 -10.480 16.375 ;
        RECT -9.070 15.335 -8.900 16.375 ;
        RECT -7.490 15.335 -7.320 16.375 ;
        RECT -5.910 15.335 -5.740 16.375 ;
        RECT -4.330 15.335 -4.160 16.375 ;
        RECT -2.750 15.335 -2.580 16.375 ;
        RECT -1.170 15.335 -1.000 16.375 ;
        RECT 0.410 15.335 0.580 16.375 ;
        RECT 1.990 15.335 2.160 16.375 ;
        RECT 3.570 15.335 3.740 16.375 ;
        RECT 5.150 15.335 5.320 16.375 ;
        RECT 6.730 15.335 6.900 16.375 ;
        RECT 8.310 15.335 8.480 16.375 ;
        RECT 9.890 15.335 10.060 16.375 ;
        RECT 11.470 15.335 11.640 16.375 ;
        RECT -20.130 13.155 -19.960 14.195 ;
        RECT -18.550 13.155 -18.380 14.195 ;
        RECT -16.970 13.155 -16.800 14.195 ;
        RECT -15.390 13.155 -15.220 14.195 ;
        RECT -13.810 13.155 -13.640 14.195 ;
        RECT -12.230 13.155 -12.060 14.195 ;
        RECT -10.650 13.155 -10.480 14.195 ;
        RECT -9.070 13.155 -8.900 14.195 ;
        RECT -7.490 13.155 -7.320 14.195 ;
        RECT -5.910 13.155 -5.740 14.195 ;
        RECT -4.330 13.155 -4.160 14.195 ;
        RECT -2.750 13.155 -2.580 14.195 ;
        RECT -1.170 13.155 -1.000 14.195 ;
        RECT 0.410 13.155 0.580 14.195 ;
        RECT 1.990 13.155 2.160 14.195 ;
        RECT 3.570 13.155 3.740 14.195 ;
        RECT 5.150 13.155 5.320 14.195 ;
        RECT 6.730 13.155 6.900 14.195 ;
        RECT 8.310 13.155 8.480 14.195 ;
        RECT 9.890 13.155 10.060 14.195 ;
        RECT 11.470 13.155 11.640 14.195 ;
        RECT -20.130 10.975 -19.960 12.015 ;
        RECT -18.550 10.975 -18.380 12.015 ;
        RECT -16.970 10.975 -16.800 12.015 ;
        RECT -15.390 10.975 -15.220 12.015 ;
        RECT -13.810 10.975 -13.640 12.015 ;
        RECT -12.230 10.975 -12.060 12.015 ;
        RECT -10.650 10.975 -10.480 12.015 ;
        RECT -9.070 10.975 -8.900 12.015 ;
        RECT -7.490 10.975 -7.320 12.015 ;
        RECT -5.910 10.975 -5.740 12.015 ;
        RECT -4.330 10.975 -4.160 12.015 ;
        RECT -2.750 10.975 -2.580 12.015 ;
        RECT -1.170 10.975 -1.000 12.015 ;
        RECT 0.410 10.975 0.580 12.015 ;
        RECT 1.990 10.975 2.160 12.015 ;
        RECT 3.570 10.975 3.740 12.015 ;
        RECT 5.150 10.975 5.320 12.015 ;
        RECT 6.730 10.975 6.900 12.015 ;
        RECT 8.310 10.975 8.480 12.015 ;
        RECT 9.890 10.975 10.060 12.015 ;
        RECT 11.470 10.975 11.640 12.015 ;
        RECT -20.130 8.795 -19.960 9.835 ;
        RECT -18.550 8.795 -18.380 9.835 ;
        RECT -16.970 8.795 -16.800 9.835 ;
        RECT -15.390 8.795 -15.220 9.835 ;
        RECT -13.810 8.795 -13.640 9.835 ;
        RECT -12.230 8.795 -12.060 9.835 ;
        RECT -10.650 8.795 -10.480 9.835 ;
        RECT -9.070 8.795 -8.900 9.835 ;
        RECT -7.490 8.795 -7.320 9.835 ;
        RECT -5.910 8.795 -5.740 9.835 ;
        RECT -4.330 8.795 -4.160 9.835 ;
        RECT -2.750 8.795 -2.580 9.835 ;
        RECT -1.170 8.795 -1.000 9.835 ;
        RECT 0.410 8.795 0.580 9.835 ;
        RECT 1.990 8.795 2.160 9.835 ;
        RECT 3.570 8.795 3.740 9.835 ;
        RECT 5.150 8.795 5.320 9.835 ;
        RECT 6.730 8.795 6.900 9.835 ;
        RECT 8.310 8.795 8.480 9.835 ;
        RECT 9.890 8.795 10.060 9.835 ;
        RECT 11.470 8.795 11.640 9.835 ;
        RECT -20.210 -5.390 -20.040 -4.350 ;
        RECT -18.630 -5.390 -18.460 -4.350 ;
        RECT -17.050 -5.390 -16.880 -4.350 ;
        RECT -15.470 -5.390 -15.300 -4.350 ;
        RECT -13.890 -5.390 -13.720 -4.350 ;
        RECT -12.310 -5.390 -12.140 -4.350 ;
        RECT -10.730 -5.390 -10.560 -4.350 ;
        RECT -9.150 -5.390 -8.980 -4.350 ;
        RECT -7.570 -5.390 -7.400 -4.350 ;
        RECT -5.990 -5.390 -5.820 -4.350 ;
        RECT -4.410 -5.390 -4.240 -4.350 ;
        RECT -2.830 -5.390 -2.660 -4.350 ;
        RECT -1.250 -5.390 -1.080 -4.350 ;
        RECT 0.330 -5.390 0.500 -4.350 ;
        RECT 1.910 -5.390 2.080 -4.350 ;
        RECT 3.490 -5.390 3.660 -4.350 ;
        RECT 5.070 -5.390 5.240 -4.350 ;
        RECT 6.650 -5.390 6.820 -4.350 ;
        RECT 8.230 -5.390 8.400 -4.350 ;
        RECT 9.810 -5.390 9.980 -4.350 ;
        RECT 11.390 -5.390 11.560 -4.350 ;
        RECT -20.210 -7.480 -20.040 -6.440 ;
        RECT -18.630 -7.480 -18.460 -6.440 ;
        RECT -17.050 -7.480 -16.880 -6.440 ;
        RECT -15.470 -7.480 -15.300 -6.440 ;
        RECT -13.890 -7.480 -13.720 -6.440 ;
        RECT -12.310 -7.480 -12.140 -6.440 ;
        RECT -10.730 -7.480 -10.560 -6.440 ;
        RECT -9.150 -7.480 -8.980 -6.440 ;
        RECT -7.570 -7.480 -7.400 -6.440 ;
        RECT -5.990 -7.480 -5.820 -6.440 ;
        RECT -4.410 -7.480 -4.240 -6.440 ;
        RECT -2.830 -7.480 -2.660 -6.440 ;
        RECT -1.250 -7.480 -1.080 -6.440 ;
        RECT 0.330 -7.480 0.500 -6.440 ;
        RECT 1.910 -7.480 2.080 -6.440 ;
        RECT 3.490 -7.480 3.660 -6.440 ;
        RECT 5.070 -7.480 5.240 -6.440 ;
        RECT 6.650 -7.480 6.820 -6.440 ;
        RECT 8.230 -7.480 8.400 -6.440 ;
        RECT 9.810 -7.480 9.980 -6.440 ;
        RECT 11.390 -7.480 11.560 -6.440 ;
        RECT -20.210 -9.570 -20.040 -8.530 ;
        RECT -18.630 -9.570 -18.460 -8.530 ;
        RECT -17.050 -9.570 -16.880 -8.530 ;
        RECT -15.470 -9.570 -15.300 -8.530 ;
        RECT -13.890 -9.570 -13.720 -8.530 ;
        RECT -12.310 -9.570 -12.140 -8.530 ;
        RECT -10.730 -9.570 -10.560 -8.530 ;
        RECT -9.150 -9.570 -8.980 -8.530 ;
        RECT -7.570 -9.570 -7.400 -8.530 ;
        RECT -5.990 -9.570 -5.820 -8.530 ;
        RECT -4.410 -9.570 -4.240 -8.530 ;
        RECT -2.830 -9.570 -2.660 -8.530 ;
        RECT -1.250 -9.570 -1.080 -8.530 ;
        RECT 0.330 -9.570 0.500 -8.530 ;
        RECT 1.910 -9.570 2.080 -8.530 ;
        RECT 3.490 -9.570 3.660 -8.530 ;
        RECT 5.070 -9.570 5.240 -8.530 ;
        RECT 6.650 -9.570 6.820 -8.530 ;
        RECT 8.230 -9.570 8.400 -8.530 ;
        RECT 9.810 -9.570 9.980 -8.530 ;
        RECT 11.390 -9.570 11.560 -8.530 ;
      LAYER met1 ;
        RECT -20.360 29.955 -19.720 30.275 ;
        RECT -18.780 29.955 -18.140 30.275 ;
        RECT -17.200 29.955 -16.560 30.275 ;
        RECT -15.620 29.955 -14.980 30.275 ;
        RECT -14.040 29.955 -13.400 30.275 ;
        RECT -12.460 29.955 -11.820 30.275 ;
        RECT -10.880 29.955 -10.240 30.275 ;
        RECT -9.300 29.955 -8.660 30.275 ;
        RECT -7.720 29.955 -7.080 30.275 ;
        RECT -6.140 29.955 -5.500 30.275 ;
        RECT -4.560 29.955 -3.920 30.275 ;
        RECT -2.980 29.955 -2.340 30.275 ;
        RECT -1.400 29.955 -0.760 30.275 ;
        RECT 0.180 29.955 0.820 30.275 ;
        RECT 1.760 29.955 2.400 30.275 ;
        RECT 3.340 29.955 3.980 30.275 ;
        RECT 4.920 29.955 5.560 30.275 ;
        RECT 6.500 29.955 7.140 30.275 ;
        RECT 8.080 29.955 8.720 30.275 ;
        RECT 9.660 29.955 10.300 30.275 ;
        RECT 11.240 29.955 11.880 30.275 ;
        RECT -20.160 29.275 -19.930 29.955 ;
        RECT -18.580 29.275 -18.350 29.955 ;
        RECT -17.000 29.275 -16.770 29.955 ;
        RECT -15.420 29.275 -15.190 29.955 ;
        RECT -13.840 29.275 -13.610 29.955 ;
        RECT -12.260 29.275 -12.030 29.955 ;
        RECT -10.680 29.275 -10.450 29.955 ;
        RECT -9.100 29.275 -8.870 29.955 ;
        RECT -7.520 29.275 -7.290 29.955 ;
        RECT -5.940 29.275 -5.710 29.955 ;
        RECT -4.360 29.275 -4.130 29.955 ;
        RECT -2.780 29.275 -2.550 29.955 ;
        RECT -1.200 29.275 -0.970 29.955 ;
        RECT 0.380 29.275 0.610 29.955 ;
        RECT 1.960 29.275 2.190 29.955 ;
        RECT 3.540 29.275 3.770 29.955 ;
        RECT 5.120 29.275 5.350 29.955 ;
        RECT 6.700 29.275 6.930 29.955 ;
        RECT 8.280 29.275 8.510 29.955 ;
        RECT 9.860 29.275 10.090 29.955 ;
        RECT 11.440 29.275 11.670 29.955 ;
        RECT -20.160 28.075 -19.930 28.095 ;
        RECT -18.580 28.075 -18.350 28.095 ;
        RECT -17.000 28.075 -16.770 28.095 ;
        RECT -15.420 28.075 -15.190 28.095 ;
        RECT -13.840 28.075 -13.610 28.095 ;
        RECT -12.260 28.075 -12.030 28.095 ;
        RECT -10.680 28.075 -10.450 28.095 ;
        RECT -9.100 28.075 -8.870 28.095 ;
        RECT -7.520 28.075 -7.290 28.095 ;
        RECT -5.940 28.075 -5.710 28.095 ;
        RECT -4.360 28.075 -4.130 28.095 ;
        RECT -2.780 28.075 -2.550 28.095 ;
        RECT -1.200 28.075 -0.970 28.095 ;
        RECT 0.380 28.075 0.610 28.095 ;
        RECT 1.960 28.075 2.190 28.095 ;
        RECT 3.540 28.075 3.770 28.095 ;
        RECT 5.120 28.075 5.350 28.095 ;
        RECT 6.700 28.075 6.930 28.095 ;
        RECT 8.280 28.075 8.510 28.095 ;
        RECT 9.860 28.075 10.090 28.095 ;
        RECT 11.440 28.075 11.670 28.095 ;
        RECT -20.360 27.755 -19.720 28.075 ;
        RECT -18.780 27.755 -18.140 28.075 ;
        RECT -17.200 27.755 -16.560 28.075 ;
        RECT -15.620 27.755 -14.980 28.075 ;
        RECT -14.040 27.755 -13.400 28.075 ;
        RECT -12.460 27.755 -11.820 28.075 ;
        RECT -10.880 27.755 -10.240 28.075 ;
        RECT -9.300 27.755 -8.660 28.075 ;
        RECT -7.720 27.755 -7.080 28.075 ;
        RECT -6.140 27.755 -5.500 28.075 ;
        RECT -4.560 27.755 -3.920 28.075 ;
        RECT -2.980 27.755 -2.340 28.075 ;
        RECT -1.400 27.755 -0.760 28.075 ;
        RECT 0.180 27.755 0.820 28.075 ;
        RECT 1.760 27.755 2.400 28.075 ;
        RECT 3.340 27.755 3.980 28.075 ;
        RECT 4.920 27.755 5.560 28.075 ;
        RECT 6.500 27.755 7.140 28.075 ;
        RECT 8.080 27.755 8.720 28.075 ;
        RECT 9.660 27.755 10.300 28.075 ;
        RECT 11.240 27.755 11.880 28.075 ;
        RECT -20.160 27.095 -19.930 27.755 ;
        RECT -18.580 27.095 -18.350 27.755 ;
        RECT -17.000 27.095 -16.770 27.755 ;
        RECT -15.420 27.095 -15.190 27.755 ;
        RECT -13.840 27.095 -13.610 27.755 ;
        RECT -12.260 27.095 -12.030 27.755 ;
        RECT -10.680 27.095 -10.450 27.755 ;
        RECT -9.100 27.095 -8.870 27.755 ;
        RECT -7.520 27.095 -7.290 27.755 ;
        RECT -5.940 27.095 -5.710 27.755 ;
        RECT -4.360 27.095 -4.130 27.755 ;
        RECT -2.780 27.095 -2.550 27.755 ;
        RECT -1.200 27.095 -0.970 27.755 ;
        RECT 0.380 27.095 0.610 27.755 ;
        RECT 1.960 27.095 2.190 27.755 ;
        RECT 3.540 27.095 3.770 27.755 ;
        RECT 5.120 27.095 5.350 27.755 ;
        RECT 6.700 27.095 6.930 27.755 ;
        RECT 8.280 27.095 8.510 27.755 ;
        RECT 9.860 27.095 10.090 27.755 ;
        RECT 11.440 27.095 11.670 27.755 ;
        RECT -20.160 25.875 -19.930 25.915 ;
        RECT -18.580 25.875 -18.350 25.915 ;
        RECT -17.000 25.875 -16.770 25.915 ;
        RECT -15.420 25.875 -15.190 25.915 ;
        RECT -13.840 25.875 -13.610 25.915 ;
        RECT -12.260 25.875 -12.030 25.915 ;
        RECT -10.680 25.875 -10.450 25.915 ;
        RECT -9.100 25.875 -8.870 25.915 ;
        RECT -7.520 25.875 -7.290 25.915 ;
        RECT -5.940 25.875 -5.710 25.915 ;
        RECT -4.360 25.875 -4.130 25.915 ;
        RECT -2.780 25.875 -2.550 25.915 ;
        RECT -1.200 25.875 -0.970 25.915 ;
        RECT 0.380 25.875 0.610 25.915 ;
        RECT 1.960 25.875 2.190 25.915 ;
        RECT 3.540 25.875 3.770 25.915 ;
        RECT 5.120 25.875 5.350 25.915 ;
        RECT 6.700 25.875 6.930 25.915 ;
        RECT 8.280 25.875 8.510 25.915 ;
        RECT 9.860 25.875 10.090 25.915 ;
        RECT 11.440 25.875 11.670 25.915 ;
        RECT -20.360 25.555 -19.720 25.875 ;
        RECT -18.780 25.555 -18.140 25.875 ;
        RECT -17.200 25.555 -16.560 25.875 ;
        RECT -15.620 25.555 -14.980 25.875 ;
        RECT -14.040 25.555 -13.400 25.875 ;
        RECT -12.460 25.555 -11.820 25.875 ;
        RECT -10.880 25.555 -10.240 25.875 ;
        RECT -9.300 25.555 -8.660 25.875 ;
        RECT -7.720 25.555 -7.080 25.875 ;
        RECT -6.140 25.555 -5.500 25.875 ;
        RECT -4.560 25.555 -3.920 25.875 ;
        RECT -2.980 25.555 -2.340 25.875 ;
        RECT -1.400 25.555 -0.760 25.875 ;
        RECT 0.180 25.555 0.820 25.875 ;
        RECT 1.760 25.555 2.400 25.875 ;
        RECT 3.340 25.555 3.980 25.875 ;
        RECT 4.920 25.555 5.560 25.875 ;
        RECT 6.500 25.555 7.140 25.875 ;
        RECT 8.080 25.555 8.720 25.875 ;
        RECT 9.660 25.555 10.300 25.875 ;
        RECT 11.240 25.555 11.880 25.875 ;
        RECT -20.160 24.915 -19.930 25.555 ;
        RECT -18.580 24.915 -18.350 25.555 ;
        RECT -17.000 24.915 -16.770 25.555 ;
        RECT -15.420 24.915 -15.190 25.555 ;
        RECT -13.840 24.915 -13.610 25.555 ;
        RECT -12.260 24.915 -12.030 25.555 ;
        RECT -10.680 24.915 -10.450 25.555 ;
        RECT -9.100 24.915 -8.870 25.555 ;
        RECT -7.520 24.915 -7.290 25.555 ;
        RECT -5.940 24.915 -5.710 25.555 ;
        RECT -4.360 24.915 -4.130 25.555 ;
        RECT -2.780 24.915 -2.550 25.555 ;
        RECT -1.200 24.915 -0.970 25.555 ;
        RECT 0.380 24.915 0.610 25.555 ;
        RECT 1.960 24.915 2.190 25.555 ;
        RECT 3.540 24.915 3.770 25.555 ;
        RECT 5.120 24.915 5.350 25.555 ;
        RECT 6.700 24.915 6.930 25.555 ;
        RECT 8.280 24.915 8.510 25.555 ;
        RECT 9.860 24.915 10.090 25.555 ;
        RECT 11.440 24.915 11.670 25.555 ;
        RECT -20.160 23.700 -19.930 23.735 ;
        RECT -18.580 23.700 -18.350 23.735 ;
        RECT -17.000 23.700 -16.770 23.735 ;
        RECT -15.420 23.700 -15.190 23.735 ;
        RECT -13.840 23.700 -13.610 23.735 ;
        RECT -12.260 23.700 -12.030 23.735 ;
        RECT -10.680 23.700 -10.450 23.735 ;
        RECT -9.100 23.700 -8.870 23.735 ;
        RECT -7.520 23.700 -7.290 23.735 ;
        RECT -5.940 23.700 -5.710 23.735 ;
        RECT -4.360 23.700 -4.130 23.735 ;
        RECT -2.780 23.700 -2.550 23.735 ;
        RECT -1.200 23.700 -0.970 23.735 ;
        RECT 0.380 23.700 0.610 23.735 ;
        RECT 1.960 23.700 2.190 23.735 ;
        RECT 3.540 23.700 3.770 23.735 ;
        RECT 5.120 23.700 5.350 23.735 ;
        RECT 6.700 23.700 6.930 23.735 ;
        RECT 8.280 23.700 8.510 23.735 ;
        RECT 9.860 23.700 10.090 23.735 ;
        RECT 11.440 23.700 11.670 23.735 ;
        RECT -20.360 23.380 -19.720 23.700 ;
        RECT -18.780 23.380 -18.140 23.700 ;
        RECT -17.200 23.380 -16.560 23.700 ;
        RECT -15.620 23.380 -14.980 23.700 ;
        RECT -14.040 23.380 -13.400 23.700 ;
        RECT -12.460 23.380 -11.820 23.700 ;
        RECT -10.880 23.380 -10.240 23.700 ;
        RECT -9.300 23.380 -8.660 23.700 ;
        RECT -7.720 23.380 -7.080 23.700 ;
        RECT -6.140 23.380 -5.500 23.700 ;
        RECT -4.560 23.380 -3.920 23.700 ;
        RECT -2.980 23.380 -2.340 23.700 ;
        RECT -1.400 23.380 -0.760 23.700 ;
        RECT 0.180 23.380 0.820 23.700 ;
        RECT 1.760 23.380 2.400 23.700 ;
        RECT 3.340 23.380 3.980 23.700 ;
        RECT 4.920 23.380 5.560 23.700 ;
        RECT 6.500 23.380 7.140 23.700 ;
        RECT 8.080 23.380 8.720 23.700 ;
        RECT 9.660 23.380 10.300 23.700 ;
        RECT 11.240 23.380 11.880 23.700 ;
        RECT -20.160 22.735 -19.930 23.380 ;
        RECT -18.580 22.735 -18.350 23.380 ;
        RECT -17.000 22.735 -16.770 23.380 ;
        RECT -15.420 22.735 -15.190 23.380 ;
        RECT -13.840 22.735 -13.610 23.380 ;
        RECT -12.260 22.735 -12.030 23.380 ;
        RECT -10.680 22.735 -10.450 23.380 ;
        RECT -9.100 22.735 -8.870 23.380 ;
        RECT -7.520 22.735 -7.290 23.380 ;
        RECT -5.940 22.735 -5.710 23.380 ;
        RECT -4.360 22.735 -4.130 23.380 ;
        RECT -2.780 22.735 -2.550 23.380 ;
        RECT -1.200 22.735 -0.970 23.380 ;
        RECT 0.380 22.735 0.610 23.380 ;
        RECT 1.960 22.735 2.190 23.380 ;
        RECT 3.540 22.735 3.770 23.380 ;
        RECT 5.120 22.735 5.350 23.380 ;
        RECT 6.700 22.735 6.930 23.380 ;
        RECT 8.280 22.735 8.510 23.380 ;
        RECT 9.860 22.735 10.090 23.380 ;
        RECT 11.440 22.735 11.670 23.380 ;
        RECT -20.360 21.255 -19.720 21.575 ;
        RECT -18.780 21.255 -18.140 21.575 ;
        RECT -17.200 21.255 -16.560 21.575 ;
        RECT -15.620 21.255 -14.980 21.575 ;
        RECT -14.040 21.255 -13.400 21.575 ;
        RECT -12.460 21.255 -11.820 21.575 ;
        RECT -10.880 21.255 -10.240 21.575 ;
        RECT -9.300 21.255 -8.660 21.575 ;
        RECT -7.720 21.255 -7.080 21.575 ;
        RECT -6.140 21.255 -5.500 21.575 ;
        RECT -4.560 21.255 -3.920 21.575 ;
        RECT -2.980 21.255 -2.340 21.575 ;
        RECT -1.400 21.255 -0.760 21.575 ;
        RECT 0.180 21.255 0.820 21.575 ;
        RECT 1.760 21.255 2.400 21.575 ;
        RECT 3.340 21.255 3.980 21.575 ;
        RECT 4.920 21.255 5.560 21.575 ;
        RECT 6.500 21.255 7.140 21.575 ;
        RECT 8.080 21.255 8.720 21.575 ;
        RECT 9.660 21.255 10.300 21.575 ;
        RECT 11.240 21.255 11.880 21.575 ;
        RECT -20.160 20.555 -19.930 21.255 ;
        RECT -18.580 20.555 -18.350 21.255 ;
        RECT -17.000 20.555 -16.770 21.255 ;
        RECT -15.420 20.555 -15.190 21.255 ;
        RECT -13.840 20.555 -13.610 21.255 ;
        RECT -12.260 20.555 -12.030 21.255 ;
        RECT -10.680 20.555 -10.450 21.255 ;
        RECT -9.100 20.555 -8.870 21.255 ;
        RECT -7.520 20.555 -7.290 21.255 ;
        RECT -5.940 20.555 -5.710 21.255 ;
        RECT -4.360 20.555 -4.130 21.255 ;
        RECT -2.780 20.555 -2.550 21.255 ;
        RECT -1.200 20.555 -0.970 21.255 ;
        RECT 0.380 20.555 0.610 21.255 ;
        RECT 1.960 20.555 2.190 21.255 ;
        RECT 3.540 20.555 3.770 21.255 ;
        RECT 5.120 20.555 5.350 21.255 ;
        RECT 6.700 20.555 6.930 21.255 ;
        RECT 8.280 20.555 8.510 21.255 ;
        RECT 9.860 20.555 10.090 21.255 ;
        RECT 11.440 20.555 11.670 21.255 ;
        RECT -20.160 18.475 -19.930 18.535 ;
        RECT -18.580 18.475 -18.350 18.535 ;
        RECT -17.000 18.475 -16.770 18.535 ;
        RECT -15.420 18.475 -15.190 18.535 ;
        RECT -13.840 18.475 -13.610 18.535 ;
        RECT -12.260 18.475 -12.030 18.535 ;
        RECT -10.680 18.475 -10.450 18.535 ;
        RECT -9.100 18.475 -8.870 18.535 ;
        RECT -7.520 18.475 -7.290 18.535 ;
        RECT -5.940 18.475 -5.710 18.535 ;
        RECT -4.360 18.475 -4.130 18.535 ;
        RECT -2.780 18.475 -2.550 18.535 ;
        RECT -1.200 18.475 -0.970 18.535 ;
        RECT 0.380 18.475 0.610 18.535 ;
        RECT 1.960 18.475 2.190 18.535 ;
        RECT 3.540 18.475 3.770 18.535 ;
        RECT 5.120 18.475 5.350 18.535 ;
        RECT 6.700 18.475 6.930 18.535 ;
        RECT 8.280 18.475 8.510 18.535 ;
        RECT 9.860 18.475 10.090 18.535 ;
        RECT 11.440 18.475 11.670 18.535 ;
        RECT -20.360 18.155 -19.720 18.475 ;
        RECT -18.780 18.155 -18.140 18.475 ;
        RECT -17.200 18.155 -16.560 18.475 ;
        RECT -15.620 18.155 -14.980 18.475 ;
        RECT -14.040 18.155 -13.400 18.475 ;
        RECT -12.460 18.155 -11.820 18.475 ;
        RECT -10.880 18.155 -10.240 18.475 ;
        RECT -9.300 18.155 -8.660 18.475 ;
        RECT -7.720 18.155 -7.080 18.475 ;
        RECT -6.140 18.155 -5.500 18.475 ;
        RECT -4.560 18.155 -3.920 18.475 ;
        RECT -2.980 18.155 -2.340 18.475 ;
        RECT -1.400 18.155 -0.760 18.475 ;
        RECT 0.180 18.155 0.820 18.475 ;
        RECT 1.760 18.155 2.400 18.475 ;
        RECT 3.340 18.155 3.980 18.475 ;
        RECT 4.920 18.155 5.560 18.475 ;
        RECT 6.500 18.155 7.140 18.475 ;
        RECT 8.080 18.155 8.720 18.475 ;
        RECT 9.660 18.155 10.300 18.475 ;
        RECT 11.240 18.155 11.880 18.475 ;
        RECT -20.160 17.535 -19.930 18.155 ;
        RECT -18.580 17.535 -18.350 18.155 ;
        RECT -17.000 17.535 -16.770 18.155 ;
        RECT -15.420 17.535 -15.190 18.155 ;
        RECT -13.840 17.535 -13.610 18.155 ;
        RECT -12.260 17.535 -12.030 18.155 ;
        RECT -10.680 17.535 -10.450 18.155 ;
        RECT -9.100 17.535 -8.870 18.155 ;
        RECT -7.520 17.535 -7.290 18.155 ;
        RECT -5.940 17.535 -5.710 18.155 ;
        RECT -4.360 17.535 -4.130 18.155 ;
        RECT -2.780 17.535 -2.550 18.155 ;
        RECT -1.200 17.535 -0.970 18.155 ;
        RECT 0.380 17.535 0.610 18.155 ;
        RECT 1.960 17.535 2.190 18.155 ;
        RECT 3.540 17.535 3.770 18.155 ;
        RECT 5.120 17.535 5.350 18.155 ;
        RECT 6.700 17.535 6.930 18.155 ;
        RECT 8.280 17.535 8.510 18.155 ;
        RECT 9.860 17.535 10.090 18.155 ;
        RECT 11.440 17.535 11.670 18.155 ;
        RECT -20.160 16.300 -19.930 16.355 ;
        RECT -18.580 16.300 -18.350 16.355 ;
        RECT -17.000 16.300 -16.770 16.355 ;
        RECT -15.420 16.300 -15.190 16.355 ;
        RECT -13.840 16.300 -13.610 16.355 ;
        RECT -12.260 16.300 -12.030 16.355 ;
        RECT -10.680 16.300 -10.450 16.355 ;
        RECT -9.100 16.300 -8.870 16.355 ;
        RECT -7.520 16.300 -7.290 16.355 ;
        RECT -5.940 16.300 -5.710 16.355 ;
        RECT -4.360 16.300 -4.130 16.355 ;
        RECT -2.780 16.300 -2.550 16.355 ;
        RECT -1.200 16.300 -0.970 16.355 ;
        RECT 0.380 16.300 0.610 16.355 ;
        RECT 1.960 16.300 2.190 16.355 ;
        RECT 3.540 16.300 3.770 16.355 ;
        RECT 5.120 16.300 5.350 16.355 ;
        RECT 6.700 16.300 6.930 16.355 ;
        RECT 8.280 16.300 8.510 16.355 ;
        RECT 9.860 16.300 10.090 16.355 ;
        RECT 11.440 16.300 11.670 16.355 ;
        RECT -20.360 15.980 -19.720 16.300 ;
        RECT -18.780 15.980 -18.140 16.300 ;
        RECT -17.200 15.980 -16.560 16.300 ;
        RECT -15.620 15.980 -14.980 16.300 ;
        RECT -14.040 15.980 -13.400 16.300 ;
        RECT -12.460 15.980 -11.820 16.300 ;
        RECT -10.880 15.980 -10.240 16.300 ;
        RECT -9.300 15.980 -8.660 16.300 ;
        RECT -7.720 15.980 -7.080 16.300 ;
        RECT -6.140 15.980 -5.500 16.300 ;
        RECT -4.560 15.980 -3.920 16.300 ;
        RECT -2.980 15.980 -2.340 16.300 ;
        RECT -1.400 15.980 -0.760 16.300 ;
        RECT 0.180 15.980 0.820 16.300 ;
        RECT 1.760 15.980 2.400 16.300 ;
        RECT 3.340 15.980 3.980 16.300 ;
        RECT 4.920 15.980 5.560 16.300 ;
        RECT 6.500 15.980 7.140 16.300 ;
        RECT 8.080 15.980 8.720 16.300 ;
        RECT 9.660 15.980 10.300 16.300 ;
        RECT 11.240 15.980 11.880 16.300 ;
        RECT -20.160 15.355 -19.930 15.980 ;
        RECT -18.580 15.355 -18.350 15.980 ;
        RECT -17.000 15.355 -16.770 15.980 ;
        RECT -15.420 15.355 -15.190 15.980 ;
        RECT -13.840 15.355 -13.610 15.980 ;
        RECT -12.260 15.355 -12.030 15.980 ;
        RECT -10.680 15.355 -10.450 15.980 ;
        RECT -9.100 15.355 -8.870 15.980 ;
        RECT -7.520 15.355 -7.290 15.980 ;
        RECT -5.940 15.355 -5.710 15.980 ;
        RECT -4.360 15.355 -4.130 15.980 ;
        RECT -2.780 15.355 -2.550 15.980 ;
        RECT -1.200 15.355 -0.970 15.980 ;
        RECT 0.380 15.355 0.610 15.980 ;
        RECT 1.960 15.355 2.190 15.980 ;
        RECT 3.540 15.355 3.770 15.980 ;
        RECT 5.120 15.355 5.350 15.980 ;
        RECT 6.700 15.355 6.930 15.980 ;
        RECT 8.280 15.355 8.510 15.980 ;
        RECT 9.860 15.355 10.090 15.980 ;
        RECT 11.440 15.355 11.670 15.980 ;
        RECT -20.160 14.125 -19.930 14.175 ;
        RECT -18.580 14.125 -18.350 14.175 ;
        RECT -17.000 14.125 -16.770 14.175 ;
        RECT -15.420 14.125 -15.190 14.175 ;
        RECT -13.840 14.125 -13.610 14.175 ;
        RECT -12.260 14.125 -12.030 14.175 ;
        RECT -10.680 14.125 -10.450 14.175 ;
        RECT -9.100 14.125 -8.870 14.175 ;
        RECT -7.520 14.125 -7.290 14.175 ;
        RECT -5.940 14.125 -5.710 14.175 ;
        RECT -4.360 14.125 -4.130 14.175 ;
        RECT -2.780 14.125 -2.550 14.175 ;
        RECT -1.200 14.125 -0.970 14.175 ;
        RECT 0.380 14.125 0.610 14.175 ;
        RECT 1.960 14.125 2.190 14.175 ;
        RECT 3.540 14.125 3.770 14.175 ;
        RECT 5.120 14.125 5.350 14.175 ;
        RECT 6.700 14.125 6.930 14.175 ;
        RECT 8.280 14.125 8.510 14.175 ;
        RECT 9.860 14.125 10.090 14.175 ;
        RECT 11.440 14.125 11.670 14.175 ;
        RECT -20.360 13.805 -19.720 14.125 ;
        RECT -18.780 13.805 -18.140 14.125 ;
        RECT -17.200 13.805 -16.560 14.125 ;
        RECT -15.620 13.805 -14.980 14.125 ;
        RECT -14.040 13.805 -13.400 14.125 ;
        RECT -12.460 13.805 -11.820 14.125 ;
        RECT -10.880 13.805 -10.240 14.125 ;
        RECT -9.300 13.805 -8.660 14.125 ;
        RECT -7.720 13.805 -7.080 14.125 ;
        RECT -6.140 13.805 -5.500 14.125 ;
        RECT -4.560 13.805 -3.920 14.125 ;
        RECT -2.980 13.805 -2.340 14.125 ;
        RECT -1.400 13.805 -0.760 14.125 ;
        RECT 0.180 13.805 0.820 14.125 ;
        RECT 1.760 13.805 2.400 14.125 ;
        RECT 3.340 13.805 3.980 14.125 ;
        RECT 4.920 13.805 5.560 14.125 ;
        RECT 6.500 13.805 7.140 14.125 ;
        RECT 8.080 13.805 8.720 14.125 ;
        RECT 9.660 13.805 10.300 14.125 ;
        RECT 11.240 13.805 11.880 14.125 ;
        RECT -20.160 13.175 -19.930 13.805 ;
        RECT -18.580 13.175 -18.350 13.805 ;
        RECT -17.000 13.175 -16.770 13.805 ;
        RECT -15.420 13.175 -15.190 13.805 ;
        RECT -13.840 13.175 -13.610 13.805 ;
        RECT -12.260 13.175 -12.030 13.805 ;
        RECT -10.680 13.175 -10.450 13.805 ;
        RECT -9.100 13.175 -8.870 13.805 ;
        RECT -7.520 13.175 -7.290 13.805 ;
        RECT -5.940 13.175 -5.710 13.805 ;
        RECT -4.360 13.175 -4.130 13.805 ;
        RECT -2.780 13.175 -2.550 13.805 ;
        RECT -1.200 13.175 -0.970 13.805 ;
        RECT 0.380 13.175 0.610 13.805 ;
        RECT 1.960 13.175 2.190 13.805 ;
        RECT 3.540 13.175 3.770 13.805 ;
        RECT 5.120 13.175 5.350 13.805 ;
        RECT 6.700 13.175 6.930 13.805 ;
        RECT 8.280 13.175 8.510 13.805 ;
        RECT 9.860 13.175 10.090 13.805 ;
        RECT 11.440 13.175 11.670 13.805 ;
        RECT -20.160 11.950 -19.930 11.995 ;
        RECT -18.580 11.950 -18.350 11.995 ;
        RECT -17.000 11.950 -16.770 11.995 ;
        RECT -15.420 11.950 -15.190 11.995 ;
        RECT -13.840 11.950 -13.610 11.995 ;
        RECT -12.260 11.950 -12.030 11.995 ;
        RECT -10.680 11.950 -10.450 11.995 ;
        RECT -9.100 11.950 -8.870 11.995 ;
        RECT -7.520 11.950 -7.290 11.995 ;
        RECT -5.940 11.950 -5.710 11.995 ;
        RECT -4.360 11.950 -4.130 11.995 ;
        RECT -2.780 11.950 -2.550 11.995 ;
        RECT -1.200 11.950 -0.970 11.995 ;
        RECT 0.380 11.950 0.610 11.995 ;
        RECT 1.960 11.950 2.190 11.995 ;
        RECT 3.540 11.950 3.770 11.995 ;
        RECT 5.120 11.950 5.350 11.995 ;
        RECT 6.700 11.950 6.930 11.995 ;
        RECT 8.280 11.950 8.510 11.995 ;
        RECT 9.860 11.950 10.090 11.995 ;
        RECT 11.440 11.950 11.670 11.995 ;
        RECT -20.360 11.630 -19.720 11.950 ;
        RECT -18.780 11.630 -18.140 11.950 ;
        RECT -17.200 11.630 -16.560 11.950 ;
        RECT -15.620 11.630 -14.980 11.950 ;
        RECT -14.040 11.630 -13.400 11.950 ;
        RECT -12.460 11.630 -11.820 11.950 ;
        RECT -10.880 11.630 -10.240 11.950 ;
        RECT -9.300 11.630 -8.660 11.950 ;
        RECT -7.720 11.630 -7.080 11.950 ;
        RECT -6.140 11.630 -5.500 11.950 ;
        RECT -4.560 11.630 -3.920 11.950 ;
        RECT -2.980 11.630 -2.340 11.950 ;
        RECT -1.400 11.630 -0.760 11.950 ;
        RECT 0.180 11.630 0.820 11.950 ;
        RECT 1.760 11.630 2.400 11.950 ;
        RECT 3.340 11.630 3.980 11.950 ;
        RECT 4.920 11.630 5.560 11.950 ;
        RECT 6.500 11.630 7.140 11.950 ;
        RECT 8.080 11.630 8.720 11.950 ;
        RECT 9.660 11.630 10.300 11.950 ;
        RECT 11.240 11.630 11.880 11.950 ;
        RECT -20.160 10.995 -19.930 11.630 ;
        RECT -18.580 10.995 -18.350 11.630 ;
        RECT -17.000 10.995 -16.770 11.630 ;
        RECT -15.420 10.995 -15.190 11.630 ;
        RECT -13.840 10.995 -13.610 11.630 ;
        RECT -12.260 10.995 -12.030 11.630 ;
        RECT -10.680 10.995 -10.450 11.630 ;
        RECT -9.100 10.995 -8.870 11.630 ;
        RECT -7.520 10.995 -7.290 11.630 ;
        RECT -5.940 10.995 -5.710 11.630 ;
        RECT -4.360 10.995 -4.130 11.630 ;
        RECT -2.780 10.995 -2.550 11.630 ;
        RECT -1.200 10.995 -0.970 11.630 ;
        RECT 0.380 10.995 0.610 11.630 ;
        RECT 1.960 10.995 2.190 11.630 ;
        RECT 3.540 10.995 3.770 11.630 ;
        RECT 5.120 10.995 5.350 11.630 ;
        RECT 6.700 10.995 6.930 11.630 ;
        RECT 8.280 10.995 8.510 11.630 ;
        RECT 9.860 10.995 10.090 11.630 ;
        RECT 11.440 10.995 11.670 11.630 ;
        RECT -20.160 9.775 -19.930 9.815 ;
        RECT -18.580 9.775 -18.350 9.815 ;
        RECT -17.000 9.775 -16.770 9.815 ;
        RECT -15.420 9.775 -15.190 9.815 ;
        RECT -13.840 9.775 -13.610 9.815 ;
        RECT -12.260 9.775 -12.030 9.815 ;
        RECT -10.680 9.775 -10.450 9.815 ;
        RECT -9.100 9.775 -8.870 9.815 ;
        RECT -7.520 9.775 -7.290 9.815 ;
        RECT -5.940 9.775 -5.710 9.815 ;
        RECT -4.360 9.775 -4.130 9.815 ;
        RECT -2.780 9.775 -2.550 9.815 ;
        RECT -1.200 9.775 -0.970 9.815 ;
        RECT 0.380 9.775 0.610 9.815 ;
        RECT 1.960 9.775 2.190 9.815 ;
        RECT 3.540 9.775 3.770 9.815 ;
        RECT 5.120 9.775 5.350 9.815 ;
        RECT 6.700 9.775 6.930 9.815 ;
        RECT 8.280 9.775 8.510 9.815 ;
        RECT 9.860 9.775 10.090 9.815 ;
        RECT 11.440 9.775 11.670 9.815 ;
        RECT -20.360 9.455 -19.720 9.775 ;
        RECT -18.780 9.455 -18.140 9.775 ;
        RECT -17.200 9.455 -16.560 9.775 ;
        RECT -15.620 9.455 -14.980 9.775 ;
        RECT -14.040 9.455 -13.400 9.775 ;
        RECT -12.460 9.455 -11.820 9.775 ;
        RECT -10.880 9.455 -10.240 9.775 ;
        RECT -9.300 9.455 -8.660 9.775 ;
        RECT -7.720 9.455 -7.080 9.775 ;
        RECT -6.140 9.455 -5.500 9.775 ;
        RECT -4.560 9.455 -3.920 9.775 ;
        RECT -2.980 9.455 -2.340 9.775 ;
        RECT -1.400 9.455 -0.760 9.775 ;
        RECT 0.180 9.455 0.820 9.775 ;
        RECT 1.760 9.455 2.400 9.775 ;
        RECT 3.340 9.455 3.980 9.775 ;
        RECT 4.920 9.455 5.560 9.775 ;
        RECT 6.500 9.455 7.140 9.775 ;
        RECT 8.080 9.455 8.720 9.775 ;
        RECT 9.660 9.455 10.300 9.775 ;
        RECT 11.240 9.455 11.880 9.775 ;
        RECT -20.160 8.815 -19.930 9.455 ;
        RECT -18.580 8.815 -18.350 9.455 ;
        RECT -17.000 8.815 -16.770 9.455 ;
        RECT -15.420 8.815 -15.190 9.455 ;
        RECT -13.840 8.815 -13.610 9.455 ;
        RECT -12.260 8.815 -12.030 9.455 ;
        RECT -10.680 8.815 -10.450 9.455 ;
        RECT -9.100 8.815 -8.870 9.455 ;
        RECT -7.520 8.815 -7.290 9.455 ;
        RECT -5.940 8.815 -5.710 9.455 ;
        RECT -4.360 8.815 -4.130 9.455 ;
        RECT -2.780 8.815 -2.550 9.455 ;
        RECT -1.200 8.815 -0.970 9.455 ;
        RECT 0.380 8.815 0.610 9.455 ;
        RECT 1.960 8.815 2.190 9.455 ;
        RECT 3.540 8.815 3.770 9.455 ;
        RECT 5.120 8.815 5.350 9.455 ;
        RECT 6.700 8.815 6.930 9.455 ;
        RECT 8.280 8.815 8.510 9.455 ;
        RECT 9.860 8.815 10.090 9.455 ;
        RECT 11.440 8.815 11.670 9.455 ;
        RECT 12.670 7.475 13.415 30.655 ;
        RECT 12.265 -0.610 13.415 5.130 ;
        RECT -20.240 -4.390 -20.010 -4.370 ;
        RECT -18.660 -4.390 -18.430 -4.370 ;
        RECT -17.080 -4.390 -16.850 -4.370 ;
        RECT -15.500 -4.390 -15.270 -4.370 ;
        RECT -13.920 -4.390 -13.690 -4.370 ;
        RECT -12.340 -4.390 -12.110 -4.370 ;
        RECT -10.760 -4.390 -10.530 -4.370 ;
        RECT -9.180 -4.390 -8.950 -4.370 ;
        RECT -7.600 -4.390 -7.370 -4.370 ;
        RECT -6.020 -4.390 -5.790 -4.370 ;
        RECT -4.440 -4.390 -4.210 -4.370 ;
        RECT -2.860 -4.390 -2.630 -4.370 ;
        RECT -1.280 -4.390 -1.050 -4.370 ;
        RECT 0.300 -4.390 0.530 -4.370 ;
        RECT 1.880 -4.390 2.110 -4.370 ;
        RECT 3.460 -4.390 3.690 -4.370 ;
        RECT 5.040 -4.390 5.270 -4.370 ;
        RECT 6.620 -4.390 6.850 -4.370 ;
        RECT 8.200 -4.390 8.430 -4.370 ;
        RECT 9.780 -4.390 10.010 -4.370 ;
        RECT 11.360 -4.390 11.590 -4.370 ;
        RECT -20.360 -4.710 -19.720 -4.390 ;
        RECT -18.780 -4.710 -18.140 -4.390 ;
        RECT -17.200 -4.710 -16.560 -4.390 ;
        RECT -15.620 -4.710 -14.980 -4.390 ;
        RECT -14.040 -4.710 -13.400 -4.390 ;
        RECT -12.460 -4.710 -11.820 -4.390 ;
        RECT -10.880 -4.710 -10.240 -4.390 ;
        RECT -9.300 -4.710 -8.660 -4.390 ;
        RECT -7.720 -4.710 -7.080 -4.390 ;
        RECT -6.140 -4.710 -5.500 -4.390 ;
        RECT -4.560 -4.710 -3.920 -4.390 ;
        RECT -2.980 -4.710 -2.340 -4.390 ;
        RECT -1.400 -4.710 -0.760 -4.390 ;
        RECT 0.180 -4.710 0.820 -4.390 ;
        RECT 1.760 -4.710 2.400 -4.390 ;
        RECT 3.340 -4.710 3.980 -4.390 ;
        RECT 4.920 -4.710 5.560 -4.390 ;
        RECT 6.500 -4.710 7.140 -4.390 ;
        RECT 8.080 -4.710 8.720 -4.390 ;
        RECT 9.660 -4.710 10.300 -4.390 ;
        RECT 11.240 -4.710 11.880 -4.390 ;
        RECT -20.240 -5.370 -20.010 -4.710 ;
        RECT -18.660 -5.370 -18.430 -4.710 ;
        RECT -17.080 -5.370 -16.850 -4.710 ;
        RECT -15.500 -5.370 -15.270 -4.710 ;
        RECT -13.920 -5.370 -13.690 -4.710 ;
        RECT -12.340 -5.370 -12.110 -4.710 ;
        RECT -10.760 -5.370 -10.530 -4.710 ;
        RECT -9.180 -5.370 -8.950 -4.710 ;
        RECT -7.600 -5.370 -7.370 -4.710 ;
        RECT -6.020 -5.370 -5.790 -4.710 ;
        RECT -4.440 -5.370 -4.210 -4.710 ;
        RECT -2.860 -5.370 -2.630 -4.710 ;
        RECT -1.280 -5.370 -1.050 -4.710 ;
        RECT 0.300 -5.370 0.530 -4.710 ;
        RECT 1.880 -5.370 2.110 -4.710 ;
        RECT 3.460 -5.370 3.690 -4.710 ;
        RECT 5.040 -5.370 5.270 -4.710 ;
        RECT 6.620 -5.370 6.850 -4.710 ;
        RECT 8.200 -5.370 8.430 -4.710 ;
        RECT 9.780 -5.370 10.010 -4.710 ;
        RECT 11.360 -5.370 11.590 -4.710 ;
        RECT -20.240 -6.480 -20.010 -6.460 ;
        RECT -18.660 -6.480 -18.430 -6.460 ;
        RECT -17.080 -6.480 -16.850 -6.460 ;
        RECT -15.500 -6.480 -15.270 -6.460 ;
        RECT -13.920 -6.480 -13.690 -6.460 ;
        RECT -12.340 -6.480 -12.110 -6.460 ;
        RECT -10.760 -6.480 -10.530 -6.460 ;
        RECT -9.180 -6.480 -8.950 -6.460 ;
        RECT -7.600 -6.480 -7.370 -6.460 ;
        RECT -6.020 -6.480 -5.790 -6.460 ;
        RECT -4.440 -6.480 -4.210 -6.460 ;
        RECT -2.860 -6.480 -2.630 -6.460 ;
        RECT -1.280 -6.480 -1.050 -6.460 ;
        RECT 0.300 -6.480 0.530 -6.460 ;
        RECT 1.880 -6.480 2.110 -6.460 ;
        RECT 3.460 -6.480 3.690 -6.460 ;
        RECT 5.040 -6.480 5.270 -6.460 ;
        RECT 6.620 -6.480 6.850 -6.460 ;
        RECT 8.200 -6.480 8.430 -6.460 ;
        RECT 9.780 -6.480 10.010 -6.460 ;
        RECT 11.360 -6.480 11.590 -6.460 ;
        RECT -20.360 -6.800 -19.720 -6.480 ;
        RECT -18.780 -6.800 -18.140 -6.480 ;
        RECT -17.200 -6.800 -16.560 -6.480 ;
        RECT -15.620 -6.800 -14.980 -6.480 ;
        RECT -14.040 -6.800 -13.400 -6.480 ;
        RECT -12.460 -6.800 -11.820 -6.480 ;
        RECT -10.880 -6.800 -10.240 -6.480 ;
        RECT -9.300 -6.800 -8.660 -6.480 ;
        RECT -7.720 -6.800 -7.080 -6.480 ;
        RECT -6.140 -6.800 -5.500 -6.480 ;
        RECT -4.560 -6.800 -3.920 -6.480 ;
        RECT -2.980 -6.800 -2.340 -6.480 ;
        RECT -1.400 -6.800 -0.760 -6.480 ;
        RECT 0.180 -6.800 0.820 -6.480 ;
        RECT 1.760 -6.800 2.400 -6.480 ;
        RECT 3.340 -6.800 3.980 -6.480 ;
        RECT 4.920 -6.800 5.560 -6.480 ;
        RECT 6.500 -6.800 7.140 -6.480 ;
        RECT 8.080 -6.800 8.720 -6.480 ;
        RECT 9.660 -6.800 10.300 -6.480 ;
        RECT 11.240 -6.800 11.880 -6.480 ;
        RECT -20.240 -7.460 -20.010 -6.800 ;
        RECT -18.660 -7.460 -18.430 -6.800 ;
        RECT -17.080 -7.460 -16.850 -6.800 ;
        RECT -15.500 -7.460 -15.270 -6.800 ;
        RECT -13.920 -7.460 -13.690 -6.800 ;
        RECT -12.340 -7.460 -12.110 -6.800 ;
        RECT -10.760 -7.460 -10.530 -6.800 ;
        RECT -9.180 -7.460 -8.950 -6.800 ;
        RECT -7.600 -7.460 -7.370 -6.800 ;
        RECT -6.020 -7.460 -5.790 -6.800 ;
        RECT -4.440 -7.460 -4.210 -6.800 ;
        RECT -2.860 -7.460 -2.630 -6.800 ;
        RECT -1.280 -7.460 -1.050 -6.800 ;
        RECT 0.300 -7.460 0.530 -6.800 ;
        RECT 1.880 -7.460 2.110 -6.800 ;
        RECT 3.460 -7.460 3.690 -6.800 ;
        RECT 5.040 -7.460 5.270 -6.800 ;
        RECT 6.620 -7.460 6.850 -6.800 ;
        RECT 8.200 -7.460 8.430 -6.800 ;
        RECT 9.780 -7.460 10.010 -6.800 ;
        RECT 11.360 -7.460 11.590 -6.800 ;
        RECT -20.240 -8.570 -20.010 -8.550 ;
        RECT -18.660 -8.570 -18.430 -8.550 ;
        RECT -17.080 -8.570 -16.850 -8.550 ;
        RECT -15.500 -8.570 -15.270 -8.550 ;
        RECT -13.920 -8.570 -13.690 -8.550 ;
        RECT -12.340 -8.570 -12.110 -8.550 ;
        RECT -10.760 -8.570 -10.530 -8.550 ;
        RECT -9.180 -8.570 -8.950 -8.550 ;
        RECT -7.600 -8.570 -7.370 -8.550 ;
        RECT -6.020 -8.570 -5.790 -8.550 ;
        RECT -4.440 -8.570 -4.210 -8.550 ;
        RECT -2.860 -8.570 -2.630 -8.550 ;
        RECT -1.280 -8.570 -1.050 -8.550 ;
        RECT 0.300 -8.570 0.530 -8.550 ;
        RECT 1.880 -8.570 2.110 -8.550 ;
        RECT 3.460 -8.570 3.690 -8.550 ;
        RECT 5.040 -8.570 5.270 -8.550 ;
        RECT 6.620 -8.570 6.850 -8.550 ;
        RECT 8.200 -8.570 8.430 -8.550 ;
        RECT 9.780 -8.570 10.010 -8.550 ;
        RECT 11.360 -8.570 11.590 -8.550 ;
        RECT -20.360 -8.890 -19.720 -8.570 ;
        RECT -18.780 -8.890 -18.140 -8.570 ;
        RECT -17.200 -8.890 -16.560 -8.570 ;
        RECT -15.620 -8.890 -14.980 -8.570 ;
        RECT -14.040 -8.890 -13.400 -8.570 ;
        RECT -12.460 -8.890 -11.820 -8.570 ;
        RECT -10.880 -8.890 -10.240 -8.570 ;
        RECT -9.300 -8.890 -8.660 -8.570 ;
        RECT -7.720 -8.890 -7.080 -8.570 ;
        RECT -6.140 -8.890 -5.500 -8.570 ;
        RECT -4.560 -8.890 -3.920 -8.570 ;
        RECT -2.980 -8.890 -2.340 -8.570 ;
        RECT -1.400 -8.890 -0.760 -8.570 ;
        RECT 0.180 -8.890 0.820 -8.570 ;
        RECT 1.760 -8.890 2.400 -8.570 ;
        RECT 3.340 -8.890 3.980 -8.570 ;
        RECT 4.920 -8.890 5.560 -8.570 ;
        RECT 6.500 -8.890 7.140 -8.570 ;
        RECT 8.080 -8.890 8.720 -8.570 ;
        RECT 9.660 -8.890 10.300 -8.570 ;
        RECT 11.240 -8.890 11.880 -8.570 ;
        RECT -20.240 -9.550 -20.010 -8.890 ;
        RECT -18.660 -9.550 -18.430 -8.890 ;
        RECT -17.080 -9.550 -16.850 -8.890 ;
        RECT -15.500 -9.550 -15.270 -8.890 ;
        RECT -13.920 -9.550 -13.690 -8.890 ;
        RECT -12.340 -9.550 -12.110 -8.890 ;
        RECT -10.760 -9.550 -10.530 -8.890 ;
        RECT -9.180 -9.550 -8.950 -8.890 ;
        RECT -7.600 -9.550 -7.370 -8.890 ;
        RECT -6.020 -9.550 -5.790 -8.890 ;
        RECT -4.440 -9.550 -4.210 -8.890 ;
        RECT -2.860 -9.550 -2.630 -8.890 ;
        RECT -1.280 -9.550 -1.050 -8.890 ;
        RECT 0.300 -9.550 0.530 -8.890 ;
        RECT 1.880 -9.550 2.110 -8.890 ;
        RECT 3.460 -9.550 3.690 -8.890 ;
        RECT 5.040 -9.550 5.270 -8.890 ;
        RECT 6.620 -9.550 6.850 -8.890 ;
        RECT 8.200 -9.550 8.430 -8.890 ;
        RECT 9.780 -9.550 10.010 -8.890 ;
        RECT 11.360 -9.550 11.590 -8.890 ;
      LAYER met2 ;
        RECT -20.405 29.955 13.415 30.650 ;
        RECT 12.265 28.450 13.415 29.955 ;
        RECT -20.405 27.755 13.415 28.450 ;
        RECT 12.265 26.250 13.415 27.755 ;
        RECT -20.405 25.555 13.415 26.250 ;
        RECT 12.265 24.075 13.415 25.555 ;
        RECT -20.405 23.380 13.415 24.075 ;
        RECT 12.265 21.950 13.415 23.380 ;
        RECT -20.405 21.255 13.415 21.950 ;
        RECT 12.265 20.010 13.415 21.255 ;
        RECT 12.350 19.870 13.415 20.010 ;
        RECT 12.265 18.850 13.415 19.870 ;
        RECT -20.405 18.155 13.415 18.850 ;
        RECT 12.265 16.675 13.415 18.155 ;
        RECT -20.405 15.980 13.415 16.675 ;
        RECT 12.265 14.500 13.415 15.980 ;
        RECT -20.405 13.805 13.415 14.500 ;
        RECT 12.265 12.325 13.415 13.805 ;
        RECT -20.405 11.630 13.415 12.325 ;
        RECT 12.265 10.150 13.415 11.630 ;
        RECT -20.405 9.455 13.415 10.150 ;
        RECT 12.265 3.165 13.415 9.455 ;
        RECT 12.265 -4.015 13.495 3.165 ;
        RECT -20.460 -4.710 13.495 -4.015 ;
        RECT 12.185 -6.105 13.495 -4.710 ;
        RECT -20.405 -6.800 13.495 -6.105 ;
        RECT 12.185 -8.195 13.495 -6.800 ;
        RECT -20.405 -8.890 13.495 -8.195 ;
    END
  END out
  PIN ena
    ANTENNAGATEAREA 0.860000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER li1 ;
        RECT 8.300 -0.095 8.800 0.075 ;
        RECT -19.340 -0.740 -18.700 -0.260 ;
        RECT 8.300 -1.645 8.800 -1.475 ;
      LAYER met1 ;
        RECT -21.805 1.625 -20.630 1.820 ;
        RECT -21.805 1.220 -18.810 1.625 ;
        RECT -21.805 0.820 -20.630 1.220 ;
        RECT -19.230 -0.230 -18.810 1.220 ;
        RECT 8.465 0.870 8.630 0.875 ;
        RECT 7.915 0.610 8.660 0.870 ;
        RECT 8.465 0.105 8.630 0.610 ;
        RECT 8.320 -0.125 8.780 0.105 ;
        RECT -19.320 -0.770 -18.720 -0.230 ;
        RECT 8.465 -1.445 8.630 -0.125 ;
        RECT 8.320 -1.675 8.780 -1.445 ;
      LAYER met2 ;
        RECT -19.145 0.660 8.660 0.870 ;
        RECT -19.145 0.075 -18.870 0.660 ;
        RECT 7.915 0.610 8.660 0.660 ;
    END
  END ena
  PIN vss
    ANTENNADIFFAREA 86.656197 ;
    PORT
      LAYER pwell ;
        RECT -25.040 -2.120 -23.030 4.710 ;
        RECT -20.010 3.585 -18.030 5.565 ;
        RECT -20.010 1.510 -18.030 3.490 ;
        RECT -16.915 1.000 1.055 1.005 ;
        RECT 4.985 1.000 9.940 1.005 ;
        RECT -20.010 -1.490 -18.030 0.490 ;
        RECT -16.915 -2.575 9.940 1.000 ;
        RECT 0.440 -2.580 5.590 -2.575 ;
        RECT -21.120 -10.840 12.470 -3.080 ;
        RECT -19.940 -17.780 11.040 -11.000 ;
      LAYER li1 ;
        RECT -20.300 5.215 -17.895 5.625 ;
        RECT -24.860 4.360 -23.210 4.530 ;
        RECT -24.860 2.340 -24.690 4.360 ;
        RECT -23.380 3.000 -23.210 4.360 ;
        RECT -20.300 3.935 -19.660 5.215 ;
        RECT -18.380 3.935 -17.895 5.215 ;
        RECT -20.300 3.140 -17.895 3.935 ;
        RECT -25.120 -1.120 -24.690 2.340 ;
        RECT -24.860 -1.770 -24.690 -1.120 ;
        RECT -24.210 -1.290 -23.860 0.870 ;
        RECT -23.410 -0.460 -23.010 3.000 ;
        RECT -20.300 1.860 -19.660 3.140 ;
        RECT -18.380 1.860 -17.895 3.140 ;
        RECT -20.300 0.985 -17.895 1.860 ;
        RECT -20.300 0.595 11.455 0.985 ;
        RECT -20.300 0.310 -16.505 0.595 ;
        RECT -20.920 0.140 -16.505 0.310 ;
        RECT -23.380 -1.770 -23.210 -0.460 ;
        RECT -20.920 -1.140 -19.655 0.140 ;
        RECT -18.380 -1.140 -16.505 0.140 ;
        RECT -20.920 -1.230 -16.505 -1.140 ;
        RECT -24.860 -1.940 -23.210 -1.770 ;
        RECT -20.915 -2.165 -16.505 -1.230 ;
        RECT -14.545 -2.165 -14.335 0.595 ;
        RECT -12.375 -2.165 -12.165 0.595 ;
        RECT -11.665 -1.305 -11.495 -0.265 ;
        RECT -10.205 -2.165 -9.995 0.595 ;
        RECT -8.035 -2.165 -7.825 0.595 ;
        RECT -5.865 -2.165 -5.655 0.595 ;
        RECT -5.155 -1.305 -4.985 -0.265 ;
        RECT -3.695 -2.165 -3.485 0.595 ;
        RECT -2.195 -1.305 -2.025 -0.265 ;
        RECT -1.525 -2.165 -1.315 0.595 ;
        RECT 0.645 0.590 5.395 0.595 ;
        RECT -0.815 -1.305 -0.645 -0.265 ;
        RECT 0.645 -2.165 0.850 0.590 ;
        RECT 1.350 -1.310 1.520 -0.270 ;
        RECT 2.930 -1.310 3.100 -0.270 ;
        RECT 4.510 -1.310 4.680 -0.270 ;
        RECT -20.915 -2.170 0.850 -2.165 ;
        RECT 5.180 -2.165 5.395 0.590 ;
        RECT 6.685 -1.305 6.855 -0.265 ;
        RECT 7.355 -2.165 7.570 0.595 ;
        RECT 9.530 0.545 11.455 0.595 ;
        RECT 9.530 -2.165 12.200 0.545 ;
        RECT 5.180 -2.170 12.200 -2.165 ;
        RECT -20.915 -2.200 12.200 -2.170 ;
        RECT -20.930 -2.590 12.200 -2.200 ;
        RECT -20.930 -3.320 12.195 -2.590 ;
        RECT -20.930 -3.400 12.230 -3.320 ;
        RECT -20.880 -3.490 12.230 -3.400 ;
        RECT -20.880 -10.430 -20.710 -3.490 ;
        RECT -19.420 -5.390 -19.250 -4.350 ;
        RECT -17.840 -5.390 -17.670 -4.350 ;
        RECT -16.260 -5.390 -16.090 -4.350 ;
        RECT -14.680 -5.390 -14.510 -4.350 ;
        RECT -13.100 -5.390 -12.930 -4.350 ;
        RECT -11.520 -5.390 -11.350 -4.350 ;
        RECT -9.940 -5.390 -9.770 -4.350 ;
        RECT -8.360 -5.390 -8.190 -4.350 ;
        RECT -6.780 -5.390 -6.610 -4.350 ;
        RECT -5.200 -5.390 -5.030 -4.350 ;
        RECT -3.620 -5.390 -3.450 -4.350 ;
        RECT -2.040 -5.390 -1.870 -4.350 ;
        RECT -0.460 -5.390 -0.290 -4.350 ;
        RECT 1.120 -5.390 1.290 -4.350 ;
        RECT 2.700 -5.390 2.870 -4.350 ;
        RECT 4.280 -5.390 4.450 -4.350 ;
        RECT 5.860 -5.390 6.030 -4.350 ;
        RECT 7.440 -5.390 7.610 -4.350 ;
        RECT 9.020 -5.390 9.190 -4.350 ;
        RECT 10.600 -5.390 10.770 -4.350 ;
        RECT -19.420 -7.480 -19.250 -6.440 ;
        RECT -17.840 -7.480 -17.670 -6.440 ;
        RECT -16.260 -7.480 -16.090 -6.440 ;
        RECT -14.680 -7.480 -14.510 -6.440 ;
        RECT -13.100 -7.480 -12.930 -6.440 ;
        RECT -11.520 -7.480 -11.350 -6.440 ;
        RECT -9.940 -7.480 -9.770 -6.440 ;
        RECT -8.360 -7.480 -8.190 -6.440 ;
        RECT -6.780 -7.480 -6.610 -6.440 ;
        RECT -5.200 -7.480 -5.030 -6.440 ;
        RECT -3.620 -7.480 -3.450 -6.440 ;
        RECT -2.040 -7.480 -1.870 -6.440 ;
        RECT -0.460 -7.480 -0.290 -6.440 ;
        RECT 1.120 -7.480 1.290 -6.440 ;
        RECT 2.700 -7.480 2.870 -6.440 ;
        RECT 4.280 -7.480 4.450 -6.440 ;
        RECT 5.860 -7.480 6.030 -6.440 ;
        RECT 7.440 -7.480 7.610 -6.440 ;
        RECT 9.020 -7.480 9.190 -6.440 ;
        RECT 10.600 -7.480 10.770 -6.440 ;
        RECT -19.420 -9.570 -19.250 -8.530 ;
        RECT -17.840 -9.570 -17.670 -8.530 ;
        RECT -16.260 -9.570 -16.090 -8.530 ;
        RECT -14.680 -9.570 -14.510 -8.530 ;
        RECT -13.100 -9.570 -12.930 -8.530 ;
        RECT -11.520 -9.570 -11.350 -8.530 ;
        RECT -9.940 -9.570 -9.770 -8.530 ;
        RECT -8.360 -9.570 -8.190 -8.530 ;
        RECT -6.780 -9.570 -6.610 -8.530 ;
        RECT -5.200 -9.570 -5.030 -8.530 ;
        RECT -3.620 -9.570 -3.450 -8.530 ;
        RECT -2.040 -9.570 -1.870 -8.530 ;
        RECT -0.460 -9.570 -0.290 -8.530 ;
        RECT 1.120 -9.570 1.290 -8.530 ;
        RECT 2.700 -9.570 2.870 -8.530 ;
        RECT 4.280 -9.570 4.450 -8.530 ;
        RECT 5.860 -9.570 6.030 -8.530 ;
        RECT 7.440 -9.570 7.610 -8.530 ;
        RECT 9.020 -9.570 9.190 -8.530 ;
        RECT 10.600 -9.570 10.770 -8.530 ;
        RECT 12.060 -10.430 12.230 -3.490 ;
        RECT -20.880 -10.600 12.230 -10.430 ;
        RECT -20.875 -11.350 12.215 -10.600 ;
        RECT -20.875 -17.430 -19.590 -11.350 ;
        RECT 10.690 -17.430 12.215 -11.350 ;
        RECT -20.875 -18.030 12.215 -17.430 ;
      LAYER met1 ;
        RECT -25.020 2.400 -24.600 2.890 ;
        RECT -23.440 2.860 -22.980 3.060 ;
        RECT -25.150 -0.070 -24.600 2.400 ;
        RECT -25.150 -1.180 -24.690 -0.070 ;
        RECT -24.220 -0.970 -23.860 0.850 ;
        RECT -23.450 -0.050 -22.980 2.860 ;
        RECT -23.440 -0.520 -22.980 -0.050 ;
        RECT -24.320 -1.740 -23.750 -0.970 ;
        RECT -21.960 -0.990 -19.900 0.170 ;
        RECT -17.685 -0.990 -16.900 0.280 ;
        RECT -5.540 -0.285 -5.065 -0.270 ;
        RECT -11.695 -0.290 -11.465 -0.285 ;
        RECT -21.960 -1.675 -16.900 -0.990 ;
        RECT -24.460 -1.860 -23.590 -1.740 ;
        RECT -21.960 -1.860 -19.900 -1.675 ;
        RECT -24.460 -2.190 -19.900 -1.860 ;
        RECT -24.310 -2.290 -19.900 -2.190 ;
        RECT -21.960 -2.730 -19.900 -2.290 ;
        RECT -17.685 -2.430 -16.900 -1.675 ;
        RECT -12.035 -1.285 -11.465 -0.290 ;
        RECT -5.540 -1.285 -4.955 -0.285 ;
        RECT -2.225 -0.295 -1.995 -0.285 ;
        RECT -0.845 -0.295 -0.615 -0.285 ;
        RECT -2.225 -1.275 -0.615 -0.295 ;
        RECT 1.320 -0.390 1.550 -0.290 ;
        RECT 2.900 -0.380 3.130 -0.290 ;
        RECT 4.480 -0.370 4.710 -0.290 ;
        RECT 6.655 -0.360 6.885 -0.285 ;
        RECT -2.225 -1.285 -1.995 -1.275 ;
        RECT -12.035 -2.655 -11.560 -1.285 ;
        RECT -5.540 -2.655 -5.065 -1.285 ;
        RECT -1.705 -2.655 -1.030 -1.275 ;
        RECT -0.845 -1.285 -0.615 -1.275 ;
        RECT 1.220 -1.310 1.630 -0.390 ;
        RECT 2.815 -1.300 3.225 -0.380 ;
        RECT 4.395 -1.290 4.805 -0.370 ;
        RECT 6.560 -1.280 6.970 -0.360 ;
        RECT 6.655 -1.285 6.885 -1.280 ;
        RECT -21.960 -2.735 -20.600 -2.730 ;
        RECT -18.535 -3.300 11.355 -2.655 ;
        RECT -19.450 -5.015 -19.220 -4.370 ;
        RECT -17.870 -5.015 -17.640 -4.370 ;
        RECT -16.290 -5.015 -16.060 -4.370 ;
        RECT -14.710 -5.015 -14.480 -4.370 ;
        RECT -13.130 -5.015 -12.900 -4.370 ;
        RECT -11.550 -5.015 -11.320 -4.370 ;
        RECT -9.970 -5.015 -9.740 -4.370 ;
        RECT -8.390 -5.015 -8.160 -4.370 ;
        RECT -6.810 -5.015 -6.580 -4.370 ;
        RECT -5.230 -5.015 -5.000 -4.370 ;
        RECT -3.650 -5.015 -3.420 -4.370 ;
        RECT -2.070 -5.015 -1.840 -4.370 ;
        RECT -0.490 -5.015 -0.260 -4.370 ;
        RECT 1.090 -5.015 1.320 -4.370 ;
        RECT 2.670 -5.015 2.900 -4.370 ;
        RECT 4.250 -5.015 4.480 -4.370 ;
        RECT 5.830 -5.015 6.060 -4.370 ;
        RECT 7.410 -5.015 7.640 -4.370 ;
        RECT 8.990 -5.015 9.220 -4.370 ;
        RECT 10.570 -5.015 10.800 -4.370 ;
        RECT -19.570 -5.335 -18.930 -5.015 ;
        RECT -17.990 -5.335 -17.350 -5.015 ;
        RECT -16.410 -5.335 -15.770 -5.015 ;
        RECT -14.830 -5.335 -14.190 -5.015 ;
        RECT -13.250 -5.335 -12.610 -5.015 ;
        RECT -11.670 -5.335 -11.030 -5.015 ;
        RECT -10.090 -5.335 -9.450 -5.015 ;
        RECT -8.510 -5.335 -7.870 -5.015 ;
        RECT -6.930 -5.335 -6.290 -5.015 ;
        RECT -5.350 -5.335 -4.710 -5.015 ;
        RECT -3.770 -5.335 -3.130 -5.015 ;
        RECT -2.190 -5.335 -1.550 -5.015 ;
        RECT -0.610 -5.335 0.030 -5.015 ;
        RECT 0.970 -5.335 1.610 -5.015 ;
        RECT 2.550 -5.335 3.190 -5.015 ;
        RECT 4.130 -5.335 4.770 -5.015 ;
        RECT 5.710 -5.335 6.350 -5.015 ;
        RECT 7.290 -5.335 7.930 -5.015 ;
        RECT 8.870 -5.335 9.510 -5.015 ;
        RECT 10.450 -5.335 11.090 -5.015 ;
        RECT -19.450 -5.370 -19.220 -5.335 ;
        RECT -17.870 -5.370 -17.640 -5.335 ;
        RECT -16.290 -5.370 -16.060 -5.335 ;
        RECT -14.710 -5.370 -14.480 -5.335 ;
        RECT -13.130 -5.370 -12.900 -5.335 ;
        RECT -11.550 -5.370 -11.320 -5.335 ;
        RECT -9.970 -5.370 -9.740 -5.335 ;
        RECT -8.390 -5.370 -8.160 -5.335 ;
        RECT -6.810 -5.370 -6.580 -5.335 ;
        RECT -5.230 -5.370 -5.000 -5.335 ;
        RECT -3.650 -5.370 -3.420 -5.335 ;
        RECT -2.070 -5.370 -1.840 -5.335 ;
        RECT -0.490 -5.370 -0.260 -5.335 ;
        RECT 1.090 -5.370 1.320 -5.335 ;
        RECT 2.670 -5.370 2.900 -5.335 ;
        RECT 4.250 -5.370 4.480 -5.335 ;
        RECT 5.830 -5.370 6.060 -5.335 ;
        RECT 7.410 -5.370 7.640 -5.335 ;
        RECT 8.990 -5.370 9.220 -5.335 ;
        RECT 10.570 -5.370 10.800 -5.335 ;
        RECT -19.450 -7.105 -19.220 -6.460 ;
        RECT -17.870 -7.105 -17.640 -6.460 ;
        RECT -16.290 -7.105 -16.060 -6.460 ;
        RECT -14.710 -7.105 -14.480 -6.460 ;
        RECT -13.130 -7.105 -12.900 -6.460 ;
        RECT -11.550 -7.105 -11.320 -6.460 ;
        RECT -9.970 -7.105 -9.740 -6.460 ;
        RECT -8.390 -7.105 -8.160 -6.460 ;
        RECT -6.810 -7.105 -6.580 -6.460 ;
        RECT -5.230 -7.105 -5.000 -6.460 ;
        RECT -3.650 -7.105 -3.420 -6.460 ;
        RECT -2.070 -7.105 -1.840 -6.460 ;
        RECT -0.490 -7.105 -0.260 -6.460 ;
        RECT 1.090 -7.105 1.320 -6.460 ;
        RECT 2.670 -7.105 2.900 -6.460 ;
        RECT 4.250 -7.105 4.480 -6.460 ;
        RECT 5.830 -7.105 6.060 -6.460 ;
        RECT 7.410 -7.105 7.640 -6.460 ;
        RECT 8.990 -7.105 9.220 -6.460 ;
        RECT 10.570 -7.105 10.800 -6.460 ;
        RECT -19.570 -7.425 -18.930 -7.105 ;
        RECT -17.990 -7.425 -17.350 -7.105 ;
        RECT -16.410 -7.425 -15.770 -7.105 ;
        RECT -14.830 -7.425 -14.190 -7.105 ;
        RECT -13.250 -7.425 -12.610 -7.105 ;
        RECT -11.670 -7.425 -11.030 -7.105 ;
        RECT -10.090 -7.425 -9.450 -7.105 ;
        RECT -8.510 -7.425 -7.870 -7.105 ;
        RECT -6.930 -7.425 -6.290 -7.105 ;
        RECT -5.350 -7.425 -4.710 -7.105 ;
        RECT -3.770 -7.425 -3.130 -7.105 ;
        RECT -2.190 -7.425 -1.550 -7.105 ;
        RECT -0.610 -7.425 0.030 -7.105 ;
        RECT 0.970 -7.425 1.610 -7.105 ;
        RECT 2.550 -7.425 3.190 -7.105 ;
        RECT 4.130 -7.425 4.770 -7.105 ;
        RECT 5.710 -7.425 6.350 -7.105 ;
        RECT 7.290 -7.425 7.930 -7.105 ;
        RECT 8.870 -7.425 9.510 -7.105 ;
        RECT 10.450 -7.425 11.090 -7.105 ;
        RECT -19.450 -7.460 -19.220 -7.425 ;
        RECT -17.870 -7.460 -17.640 -7.425 ;
        RECT -16.290 -7.460 -16.060 -7.425 ;
        RECT -14.710 -7.460 -14.480 -7.425 ;
        RECT -13.130 -7.460 -12.900 -7.425 ;
        RECT -11.550 -7.460 -11.320 -7.425 ;
        RECT -9.970 -7.460 -9.740 -7.425 ;
        RECT -8.390 -7.460 -8.160 -7.425 ;
        RECT -6.810 -7.460 -6.580 -7.425 ;
        RECT -5.230 -7.460 -5.000 -7.425 ;
        RECT -3.650 -7.460 -3.420 -7.425 ;
        RECT -2.070 -7.460 -1.840 -7.425 ;
        RECT -0.490 -7.460 -0.260 -7.425 ;
        RECT 1.090 -7.460 1.320 -7.425 ;
        RECT 2.670 -7.460 2.900 -7.425 ;
        RECT 4.250 -7.460 4.480 -7.425 ;
        RECT 5.830 -7.460 6.060 -7.425 ;
        RECT 7.410 -7.460 7.640 -7.425 ;
        RECT 8.990 -7.460 9.220 -7.425 ;
        RECT 10.570 -7.460 10.800 -7.425 ;
        RECT -19.450 -9.195 -19.220 -8.550 ;
        RECT -17.870 -9.195 -17.640 -8.550 ;
        RECT -16.290 -9.195 -16.060 -8.550 ;
        RECT -14.710 -9.195 -14.480 -8.550 ;
        RECT -13.130 -9.195 -12.900 -8.550 ;
        RECT -11.550 -9.195 -11.320 -8.550 ;
        RECT -9.970 -9.195 -9.740 -8.550 ;
        RECT -8.390 -9.195 -8.160 -8.550 ;
        RECT -6.810 -9.195 -6.580 -8.550 ;
        RECT -5.230 -9.195 -5.000 -8.550 ;
        RECT -3.650 -9.195 -3.420 -8.550 ;
        RECT -2.070 -9.195 -1.840 -8.550 ;
        RECT -0.490 -9.195 -0.260 -8.550 ;
        RECT 1.090 -9.195 1.320 -8.550 ;
        RECT 2.670 -9.195 2.900 -8.550 ;
        RECT 4.250 -9.195 4.480 -8.550 ;
        RECT 5.830 -9.195 6.060 -8.550 ;
        RECT 7.410 -9.195 7.640 -8.550 ;
        RECT 8.990 -9.195 9.220 -8.550 ;
        RECT 10.570 -9.195 10.800 -8.550 ;
        RECT -19.570 -9.515 -18.930 -9.195 ;
        RECT -17.990 -9.515 -17.350 -9.195 ;
        RECT -16.410 -9.515 -15.770 -9.195 ;
        RECT -14.830 -9.515 -14.190 -9.195 ;
        RECT -13.250 -9.515 -12.610 -9.195 ;
        RECT -11.670 -9.515 -11.030 -9.195 ;
        RECT -10.090 -9.515 -9.450 -9.195 ;
        RECT -8.510 -9.515 -7.870 -9.195 ;
        RECT -6.930 -9.515 -6.290 -9.195 ;
        RECT -5.350 -9.515 -4.710 -9.195 ;
        RECT -3.770 -9.515 -3.130 -9.195 ;
        RECT -2.190 -9.515 -1.550 -9.195 ;
        RECT -0.610 -9.515 0.030 -9.195 ;
        RECT 0.970 -9.515 1.610 -9.195 ;
        RECT 2.550 -9.515 3.190 -9.195 ;
        RECT 4.130 -9.515 4.770 -9.195 ;
        RECT 5.710 -9.515 6.350 -9.195 ;
        RECT 7.290 -9.515 7.930 -9.195 ;
        RECT 8.870 -9.515 9.510 -9.195 ;
        RECT 10.450 -9.515 11.090 -9.195 ;
        RECT -19.450 -9.550 -19.220 -9.515 ;
        RECT -17.870 -9.550 -17.640 -9.515 ;
        RECT -16.290 -9.550 -16.060 -9.515 ;
        RECT -14.710 -9.550 -14.480 -9.515 ;
        RECT -13.130 -9.550 -12.900 -9.515 ;
        RECT -11.550 -9.550 -11.320 -9.515 ;
        RECT -9.970 -9.550 -9.740 -9.515 ;
        RECT -8.390 -9.550 -8.160 -9.515 ;
        RECT -6.810 -9.550 -6.580 -9.515 ;
        RECT -5.230 -9.550 -5.000 -9.515 ;
        RECT -3.650 -9.550 -3.420 -9.515 ;
        RECT -2.070 -9.550 -1.840 -9.515 ;
        RECT -0.490 -9.550 -0.260 -9.515 ;
        RECT 1.090 -9.550 1.320 -9.515 ;
        RECT 2.670 -9.550 2.900 -9.515 ;
        RECT 4.250 -9.550 4.480 -9.515 ;
        RECT 5.830 -9.550 6.060 -9.515 ;
        RECT 7.410 -9.550 7.640 -9.515 ;
        RECT 8.990 -9.550 9.220 -9.515 ;
        RECT 10.570 -9.550 10.800 -9.515 ;
        RECT -21.960 -11.275 11.765 -10.495 ;
        RECT -21.960 -12.360 -19.970 -11.275 ;
        RECT -20.625 -17.585 -19.970 -12.360 ;
        RECT -16.265 -16.860 -15.265 -11.275 ;
        RECT -14.265 -17.585 -13.265 -12.130 ;
        RECT -12.265 -16.860 -11.265 -11.275 ;
        RECT -10.265 -17.585 -9.265 -12.130 ;
        RECT -8.265 -16.860 -7.265 -11.275 ;
        RECT -6.265 -17.585 -5.265 -12.130 ;
        RECT -4.265 -16.860 -3.265 -11.275 ;
        RECT -2.265 -17.585 -1.265 -12.130 ;
        RECT -0.265 -16.860 0.735 -11.275 ;
        RECT 1.735 -17.585 2.735 -12.130 ;
        RECT 3.735 -16.860 4.735 -11.275 ;
        RECT 5.735 -17.585 6.735 -12.130 ;
        RECT 11.450 -17.585 12.010 -12.390 ;
        RECT -20.625 -18.030 12.010 -17.585 ;
      LAYER met2 ;
        RECT -25.170 2.940 -24.660 4.310 ;
        RECT -25.170 -0.120 -24.650 2.940 ;
        RECT -31.350 -1.890 -29.710 -1.650 ;
        RECT -25.170 -1.740 -24.660 -0.120 ;
        RECT -24.410 -1.740 -23.640 -1.690 ;
        RECT -23.400 -1.740 -22.710 4.310 ;
        RECT -21.960 -1.740 -20.605 0.220 ;
        RECT -31.350 -1.900 -25.540 -1.890 ;
        RECT -25.170 -1.900 -20.605 -1.740 ;
        RECT -31.350 -2.655 -20.605 -1.900 ;
        RECT 1.195 -2.655 1.630 -0.395 ;
        RECT 2.800 -2.655 3.235 -0.360 ;
        RECT 4.395 -2.655 4.830 -0.360 ;
        RECT 6.560 -2.655 6.995 -0.365 ;
        RECT -31.350 -2.900 11.355 -2.655 ;
        RECT -31.350 -2.910 -25.540 -2.900 ;
        RECT -23.400 -2.910 -22.710 -2.900 ;
        RECT -31.350 -3.200 -29.710 -2.910 ;
        RECT -29.020 -2.920 -27.810 -2.910 ;
        RECT -21.960 -3.425 11.355 -2.900 ;
        RECT -21.960 -5.015 -20.605 -3.425 ;
        RECT -21.965 -5.710 11.915 -5.015 ;
        RECT -21.960 -7.105 -20.605 -5.710 ;
        RECT -21.960 -7.800 11.915 -7.105 ;
        RECT -21.960 -9.195 -20.605 -7.800 ;
        RECT -21.960 -9.890 11.915 -9.195 ;
        RECT -21.960 -12.360 -20.605 -9.890 ;
      LAYER met3 ;
        RECT -31.250 -3.065 -29.800 -1.725 ;
      LAYER met4 ;
        RECT -31.330 36.050 21.520 37.910 ;
        RECT -31.205 -3.055 -29.845 -1.745 ;
        RECT -31.330 -24.580 21.550 -22.730 ;
      LAYER met5 ;
        RECT -31.330 35.580 -29.720 37.910 ;
        RECT -31.340 -21.200 -29.720 35.580 ;
        RECT -31.330 -24.570 -29.720 -21.200 ;
        RECT 19.910 -22.730 21.520 37.920 ;
        RECT 19.910 -24.580 21.560 -22.730 ;
    END
  END vss
  PIN inp
    ANTENNAGATEAREA 2.360000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER li1 ;
        RECT -19.340 4.335 -18.700 4.815 ;
        RECT -24.210 1.720 -23.860 3.880 ;
        RECT -3.480 2.795 -2.980 2.965 ;
        RECT -2.690 2.795 -2.190 2.965 ;
        RECT -13.605 -0.095 -13.105 0.075 ;
        RECT -7.095 -0.095 -6.595 0.075 ;
        RECT -13.605 -1.645 -13.105 -1.475 ;
        RECT -7.095 -1.645 -6.595 -1.475 ;
      LAYER met1 ;
        RECT -21.805 4.845 -19.040 5.095 ;
        RECT -21.805 4.750 -18.720 4.845 ;
        RECT -24.310 4.305 -18.720 4.750 ;
        RECT -24.310 4.290 -19.040 4.305 ;
        RECT -24.290 3.610 -23.720 4.290 ;
        RECT -21.805 4.095 -19.040 4.290 ;
        RECT -24.190 1.700 -23.830 3.610 ;
        RECT -3.460 2.765 -3.000 2.995 ;
        RECT -2.670 2.765 -2.210 2.995 ;
        RECT -3.325 1.875 -3.120 2.765 ;
        RECT -2.510 1.875 -2.305 2.765 ;
        RECT -13.975 1.615 -13.210 1.875 ;
        RECT -7.475 1.615 -6.710 1.875 ;
        RECT -3.325 1.615 -2.305 1.875 ;
        RECT -13.465 0.105 -13.265 1.615 ;
        RECT -6.945 0.105 -6.750 1.615 ;
        RECT -13.585 -0.125 -13.125 0.105 ;
        RECT -7.075 -0.125 -6.615 0.105 ;
        RECT -13.465 -1.445 -13.265 -0.125 ;
        RECT -6.945 -1.445 -6.750 -0.125 ;
        RECT -13.585 -1.675 -13.125 -1.445 ;
        RECT -7.075 -1.675 -6.615 -1.445 ;
      LAYER met2 ;
        RECT -20.720 4.370 -19.040 5.095 ;
        RECT -20.720 4.095 -17.565 4.370 ;
        RECT -17.840 1.865 -17.565 4.095 ;
        RECT -13.975 1.865 -13.210 1.875 ;
        RECT -7.475 1.865 -6.710 1.875 ;
        RECT -3.325 1.865 -2.305 1.875 ;
        RECT -17.840 1.615 -2.305 1.865 ;
    END
  END inp
  PIN inm
    ANTENNAGATEAREA 2.360000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER li1 ;
        RECT -0.560 2.795 -0.060 2.965 ;
        RECT 0.230 2.795 0.730 2.965 ;
        RECT -19.340 2.260 -18.700 2.740 ;
        RECT -15.775 -0.095 -15.275 0.075 ;
        RECT -9.265 -0.095 -8.765 0.075 ;
        RECT -15.775 -1.645 -15.275 -1.475 ;
        RECT -9.265 -1.645 -8.765 -1.475 ;
      LAYER met1 ;
        RECT -21.805 2.770 -18.810 3.445 ;
        RECT -21.805 2.445 -18.720 2.770 ;
        RECT -0.540 2.765 -0.080 2.995 ;
        RECT 0.250 2.765 0.710 2.995 ;
        RECT -19.320 2.230 -18.720 2.445 ;
        RECT -0.425 1.395 -0.220 2.765 ;
        RECT 0.370 1.395 0.575 2.765 ;
        RECT -16.140 1.135 -15.375 1.395 ;
        RECT -9.635 1.135 -8.870 1.395 ;
        RECT -0.430 1.135 0.580 1.395 ;
        RECT -15.615 0.105 -15.420 1.135 ;
        RECT -9.110 0.105 -8.905 1.135 ;
        RECT -15.755 -0.125 -15.295 0.105 ;
        RECT -9.245 -0.125 -8.785 0.105 ;
        RECT -15.615 -1.445 -15.420 -0.125 ;
        RECT -9.110 -1.445 -8.905 -0.125 ;
        RECT -15.755 -1.675 -15.295 -1.445 ;
        RECT -9.245 -1.675 -8.785 -1.445 ;
      LAYER met2 ;
        RECT -20.720 2.445 -18.810 3.445 ;
        RECT -19.130 1.385 -18.810 2.445 ;
        RECT -16.140 1.385 -15.375 1.395 ;
        RECT -9.635 1.385 -8.870 1.395 ;
        RECT -0.445 1.385 0.590 1.395 ;
        RECT -19.130 1.135 0.590 1.385 ;
        RECT -0.445 1.120 0.590 1.135 ;
    END
  END inm
  OBS
      LAYER li1 ;
        RECT -19.900 30.510 -19.400 30.680 ;
        RECT -19.110 30.510 -18.610 30.680 ;
        RECT -18.320 30.510 -17.820 30.680 ;
        RECT -17.530 30.510 -17.030 30.680 ;
        RECT -16.740 30.510 -16.240 30.680 ;
        RECT -15.950 30.510 -15.450 30.680 ;
        RECT -15.160 30.510 -14.660 30.680 ;
        RECT -14.370 30.510 -13.870 30.680 ;
        RECT -13.580 30.510 -13.080 30.680 ;
        RECT -12.790 30.510 -12.290 30.680 ;
        RECT -12.000 30.510 -11.500 30.680 ;
        RECT -11.210 30.510 -10.710 30.680 ;
        RECT -10.420 30.510 -9.920 30.680 ;
        RECT -9.630 30.510 -9.130 30.680 ;
        RECT -8.840 30.510 -8.340 30.680 ;
        RECT -8.050 30.510 -7.550 30.680 ;
        RECT -7.260 30.510 -6.760 30.680 ;
        RECT -6.470 30.510 -5.970 30.680 ;
        RECT -5.680 30.510 -5.180 30.680 ;
        RECT -4.890 30.510 -4.390 30.680 ;
        RECT -4.100 30.510 -3.600 30.680 ;
        RECT -3.310 30.510 -2.810 30.680 ;
        RECT -2.520 30.510 -2.020 30.680 ;
        RECT -1.730 30.510 -1.230 30.680 ;
        RECT -0.940 30.510 -0.440 30.680 ;
        RECT -0.150 30.510 0.350 30.680 ;
        RECT 0.640 30.510 1.140 30.680 ;
        RECT 1.430 30.510 1.930 30.680 ;
        RECT 2.220 30.510 2.720 30.680 ;
        RECT 3.010 30.510 3.510 30.680 ;
        RECT 3.800 30.510 4.300 30.680 ;
        RECT 4.590 30.510 5.090 30.680 ;
        RECT 5.380 30.510 5.880 30.680 ;
        RECT 6.170 30.510 6.670 30.680 ;
        RECT 6.960 30.510 7.460 30.680 ;
        RECT 7.750 30.510 8.250 30.680 ;
        RECT 8.540 30.510 9.040 30.680 ;
        RECT 9.330 30.510 9.830 30.680 ;
        RECT 10.120 30.510 10.620 30.680 ;
        RECT 10.910 30.510 11.410 30.680 ;
        RECT -19.900 28.870 -19.400 29.040 ;
        RECT -19.110 28.870 -18.610 29.040 ;
        RECT -18.320 28.870 -17.820 29.040 ;
        RECT -17.530 28.870 -17.030 29.040 ;
        RECT -16.740 28.870 -16.240 29.040 ;
        RECT -15.950 28.870 -15.450 29.040 ;
        RECT -15.160 28.870 -14.660 29.040 ;
        RECT -14.370 28.870 -13.870 29.040 ;
        RECT -13.580 28.870 -13.080 29.040 ;
        RECT -12.790 28.870 -12.290 29.040 ;
        RECT -12.000 28.870 -11.500 29.040 ;
        RECT -11.210 28.870 -10.710 29.040 ;
        RECT -10.420 28.870 -9.920 29.040 ;
        RECT -9.630 28.870 -9.130 29.040 ;
        RECT -8.840 28.870 -8.340 29.040 ;
        RECT -8.050 28.870 -7.550 29.040 ;
        RECT -7.260 28.870 -6.760 29.040 ;
        RECT -6.470 28.870 -5.970 29.040 ;
        RECT -5.680 28.870 -5.180 29.040 ;
        RECT -4.890 28.870 -4.390 29.040 ;
        RECT -4.100 28.870 -3.600 29.040 ;
        RECT -3.310 28.870 -2.810 29.040 ;
        RECT -2.520 28.870 -2.020 29.040 ;
        RECT -1.730 28.870 -1.230 29.040 ;
        RECT -0.940 28.870 -0.440 29.040 ;
        RECT -0.150 28.870 0.350 29.040 ;
        RECT 0.640 28.870 1.140 29.040 ;
        RECT 1.430 28.870 1.930 29.040 ;
        RECT 2.220 28.870 2.720 29.040 ;
        RECT 3.010 28.870 3.510 29.040 ;
        RECT 3.800 28.870 4.300 29.040 ;
        RECT 4.590 28.870 5.090 29.040 ;
        RECT 5.380 28.870 5.880 29.040 ;
        RECT 6.170 28.870 6.670 29.040 ;
        RECT 6.960 28.870 7.460 29.040 ;
        RECT 7.750 28.870 8.250 29.040 ;
        RECT 8.540 28.870 9.040 29.040 ;
        RECT 9.330 28.870 9.830 29.040 ;
        RECT 10.120 28.870 10.620 29.040 ;
        RECT 10.910 28.870 11.410 29.040 ;
        RECT -19.900 28.330 -19.400 28.500 ;
        RECT -19.110 28.330 -18.610 28.500 ;
        RECT -18.320 28.330 -17.820 28.500 ;
        RECT -17.530 28.330 -17.030 28.500 ;
        RECT -16.740 28.330 -16.240 28.500 ;
        RECT -15.950 28.330 -15.450 28.500 ;
        RECT -15.160 28.330 -14.660 28.500 ;
        RECT -14.370 28.330 -13.870 28.500 ;
        RECT -13.580 28.330 -13.080 28.500 ;
        RECT -12.790 28.330 -12.290 28.500 ;
        RECT -12.000 28.330 -11.500 28.500 ;
        RECT -11.210 28.330 -10.710 28.500 ;
        RECT -10.420 28.330 -9.920 28.500 ;
        RECT -9.630 28.330 -9.130 28.500 ;
        RECT -8.840 28.330 -8.340 28.500 ;
        RECT -8.050 28.330 -7.550 28.500 ;
        RECT -7.260 28.330 -6.760 28.500 ;
        RECT -6.470 28.330 -5.970 28.500 ;
        RECT -5.680 28.330 -5.180 28.500 ;
        RECT -4.890 28.330 -4.390 28.500 ;
        RECT -4.100 28.330 -3.600 28.500 ;
        RECT -3.310 28.330 -2.810 28.500 ;
        RECT -2.520 28.330 -2.020 28.500 ;
        RECT -1.730 28.330 -1.230 28.500 ;
        RECT -0.940 28.330 -0.440 28.500 ;
        RECT -0.150 28.330 0.350 28.500 ;
        RECT 0.640 28.330 1.140 28.500 ;
        RECT 1.430 28.330 1.930 28.500 ;
        RECT 2.220 28.330 2.720 28.500 ;
        RECT 3.010 28.330 3.510 28.500 ;
        RECT 3.800 28.330 4.300 28.500 ;
        RECT 4.590 28.330 5.090 28.500 ;
        RECT 5.380 28.330 5.880 28.500 ;
        RECT 6.170 28.330 6.670 28.500 ;
        RECT 6.960 28.330 7.460 28.500 ;
        RECT 7.750 28.330 8.250 28.500 ;
        RECT 8.540 28.330 9.040 28.500 ;
        RECT 9.330 28.330 9.830 28.500 ;
        RECT 10.120 28.330 10.620 28.500 ;
        RECT 10.910 28.330 11.410 28.500 ;
        RECT -19.900 26.690 -19.400 26.860 ;
        RECT -19.110 26.690 -18.610 26.860 ;
        RECT -18.320 26.690 -17.820 26.860 ;
        RECT -17.530 26.690 -17.030 26.860 ;
        RECT -16.740 26.690 -16.240 26.860 ;
        RECT -15.950 26.690 -15.450 26.860 ;
        RECT -15.160 26.690 -14.660 26.860 ;
        RECT -14.370 26.690 -13.870 26.860 ;
        RECT -13.580 26.690 -13.080 26.860 ;
        RECT -12.790 26.690 -12.290 26.860 ;
        RECT -12.000 26.690 -11.500 26.860 ;
        RECT -11.210 26.690 -10.710 26.860 ;
        RECT -10.420 26.690 -9.920 26.860 ;
        RECT -9.630 26.690 -9.130 26.860 ;
        RECT -8.840 26.690 -8.340 26.860 ;
        RECT -8.050 26.690 -7.550 26.860 ;
        RECT -7.260 26.690 -6.760 26.860 ;
        RECT -6.470 26.690 -5.970 26.860 ;
        RECT -5.680 26.690 -5.180 26.860 ;
        RECT -4.890 26.690 -4.390 26.860 ;
        RECT -4.100 26.690 -3.600 26.860 ;
        RECT -3.310 26.690 -2.810 26.860 ;
        RECT -2.520 26.690 -2.020 26.860 ;
        RECT -1.730 26.690 -1.230 26.860 ;
        RECT -0.940 26.690 -0.440 26.860 ;
        RECT -0.150 26.690 0.350 26.860 ;
        RECT 0.640 26.690 1.140 26.860 ;
        RECT 1.430 26.690 1.930 26.860 ;
        RECT 2.220 26.690 2.720 26.860 ;
        RECT 3.010 26.690 3.510 26.860 ;
        RECT 3.800 26.690 4.300 26.860 ;
        RECT 4.590 26.690 5.090 26.860 ;
        RECT 5.380 26.690 5.880 26.860 ;
        RECT 6.170 26.690 6.670 26.860 ;
        RECT 6.960 26.690 7.460 26.860 ;
        RECT 7.750 26.690 8.250 26.860 ;
        RECT 8.540 26.690 9.040 26.860 ;
        RECT 9.330 26.690 9.830 26.860 ;
        RECT 10.120 26.690 10.620 26.860 ;
        RECT 10.910 26.690 11.410 26.860 ;
        RECT -19.900 26.150 -19.400 26.320 ;
        RECT -19.110 26.150 -18.610 26.320 ;
        RECT -18.320 26.150 -17.820 26.320 ;
        RECT -17.530 26.150 -17.030 26.320 ;
        RECT -16.740 26.150 -16.240 26.320 ;
        RECT -15.950 26.150 -15.450 26.320 ;
        RECT -15.160 26.150 -14.660 26.320 ;
        RECT -14.370 26.150 -13.870 26.320 ;
        RECT -13.580 26.150 -13.080 26.320 ;
        RECT -12.790 26.150 -12.290 26.320 ;
        RECT -12.000 26.150 -11.500 26.320 ;
        RECT -11.210 26.150 -10.710 26.320 ;
        RECT -10.420 26.150 -9.920 26.320 ;
        RECT -9.630 26.150 -9.130 26.320 ;
        RECT -8.840 26.150 -8.340 26.320 ;
        RECT -8.050 26.150 -7.550 26.320 ;
        RECT -7.260 26.150 -6.760 26.320 ;
        RECT -6.470 26.150 -5.970 26.320 ;
        RECT -5.680 26.150 -5.180 26.320 ;
        RECT -4.890 26.150 -4.390 26.320 ;
        RECT -4.100 26.150 -3.600 26.320 ;
        RECT -3.310 26.150 -2.810 26.320 ;
        RECT -2.520 26.150 -2.020 26.320 ;
        RECT -1.730 26.150 -1.230 26.320 ;
        RECT -0.940 26.150 -0.440 26.320 ;
        RECT -0.150 26.150 0.350 26.320 ;
        RECT 0.640 26.150 1.140 26.320 ;
        RECT 1.430 26.150 1.930 26.320 ;
        RECT 2.220 26.150 2.720 26.320 ;
        RECT 3.010 26.150 3.510 26.320 ;
        RECT 3.800 26.150 4.300 26.320 ;
        RECT 4.590 26.150 5.090 26.320 ;
        RECT 5.380 26.150 5.880 26.320 ;
        RECT 6.170 26.150 6.670 26.320 ;
        RECT 6.960 26.150 7.460 26.320 ;
        RECT 7.750 26.150 8.250 26.320 ;
        RECT 8.540 26.150 9.040 26.320 ;
        RECT 9.330 26.150 9.830 26.320 ;
        RECT 10.120 26.150 10.620 26.320 ;
        RECT 10.910 26.150 11.410 26.320 ;
        RECT -19.900 24.510 -19.400 24.680 ;
        RECT -19.110 24.510 -18.610 24.680 ;
        RECT -18.320 24.510 -17.820 24.680 ;
        RECT -17.530 24.510 -17.030 24.680 ;
        RECT -16.740 24.510 -16.240 24.680 ;
        RECT -15.950 24.510 -15.450 24.680 ;
        RECT -15.160 24.510 -14.660 24.680 ;
        RECT -14.370 24.510 -13.870 24.680 ;
        RECT -13.580 24.510 -13.080 24.680 ;
        RECT -12.790 24.510 -12.290 24.680 ;
        RECT -12.000 24.510 -11.500 24.680 ;
        RECT -11.210 24.510 -10.710 24.680 ;
        RECT -10.420 24.510 -9.920 24.680 ;
        RECT -9.630 24.510 -9.130 24.680 ;
        RECT -8.840 24.510 -8.340 24.680 ;
        RECT -8.050 24.510 -7.550 24.680 ;
        RECT -7.260 24.510 -6.760 24.680 ;
        RECT -6.470 24.510 -5.970 24.680 ;
        RECT -5.680 24.510 -5.180 24.680 ;
        RECT -4.890 24.510 -4.390 24.680 ;
        RECT -4.100 24.510 -3.600 24.680 ;
        RECT -3.310 24.510 -2.810 24.680 ;
        RECT -2.520 24.510 -2.020 24.680 ;
        RECT -1.730 24.510 -1.230 24.680 ;
        RECT -0.940 24.510 -0.440 24.680 ;
        RECT -0.150 24.510 0.350 24.680 ;
        RECT 0.640 24.510 1.140 24.680 ;
        RECT 1.430 24.510 1.930 24.680 ;
        RECT 2.220 24.510 2.720 24.680 ;
        RECT 3.010 24.510 3.510 24.680 ;
        RECT 3.800 24.510 4.300 24.680 ;
        RECT 4.590 24.510 5.090 24.680 ;
        RECT 5.380 24.510 5.880 24.680 ;
        RECT 6.170 24.510 6.670 24.680 ;
        RECT 6.960 24.510 7.460 24.680 ;
        RECT 7.750 24.510 8.250 24.680 ;
        RECT 8.540 24.510 9.040 24.680 ;
        RECT 9.330 24.510 9.830 24.680 ;
        RECT 10.120 24.510 10.620 24.680 ;
        RECT 10.910 24.510 11.410 24.680 ;
        RECT -19.900 23.970 -19.400 24.140 ;
        RECT -19.110 23.970 -18.610 24.140 ;
        RECT -18.320 23.970 -17.820 24.140 ;
        RECT -17.530 23.970 -17.030 24.140 ;
        RECT -16.740 23.970 -16.240 24.140 ;
        RECT -15.950 23.970 -15.450 24.140 ;
        RECT -15.160 23.970 -14.660 24.140 ;
        RECT -14.370 23.970 -13.870 24.140 ;
        RECT -13.580 23.970 -13.080 24.140 ;
        RECT -12.790 23.970 -12.290 24.140 ;
        RECT -12.000 23.970 -11.500 24.140 ;
        RECT -11.210 23.970 -10.710 24.140 ;
        RECT -10.420 23.970 -9.920 24.140 ;
        RECT -9.630 23.970 -9.130 24.140 ;
        RECT -8.840 23.970 -8.340 24.140 ;
        RECT -8.050 23.970 -7.550 24.140 ;
        RECT -7.260 23.970 -6.760 24.140 ;
        RECT -6.470 23.970 -5.970 24.140 ;
        RECT -5.680 23.970 -5.180 24.140 ;
        RECT -4.890 23.970 -4.390 24.140 ;
        RECT -4.100 23.970 -3.600 24.140 ;
        RECT -3.310 23.970 -2.810 24.140 ;
        RECT -2.520 23.970 -2.020 24.140 ;
        RECT -1.730 23.970 -1.230 24.140 ;
        RECT -0.940 23.970 -0.440 24.140 ;
        RECT -0.150 23.970 0.350 24.140 ;
        RECT 0.640 23.970 1.140 24.140 ;
        RECT 1.430 23.970 1.930 24.140 ;
        RECT 2.220 23.970 2.720 24.140 ;
        RECT 3.010 23.970 3.510 24.140 ;
        RECT 3.800 23.970 4.300 24.140 ;
        RECT 4.590 23.970 5.090 24.140 ;
        RECT 5.380 23.970 5.880 24.140 ;
        RECT 6.170 23.970 6.670 24.140 ;
        RECT 6.960 23.970 7.460 24.140 ;
        RECT 7.750 23.970 8.250 24.140 ;
        RECT 8.540 23.970 9.040 24.140 ;
        RECT 9.330 23.970 9.830 24.140 ;
        RECT 10.120 23.970 10.620 24.140 ;
        RECT 10.910 23.970 11.410 24.140 ;
        RECT -19.900 22.330 -19.400 22.500 ;
        RECT -19.110 22.330 -18.610 22.500 ;
        RECT -18.320 22.330 -17.820 22.500 ;
        RECT -17.530 22.330 -17.030 22.500 ;
        RECT -16.740 22.330 -16.240 22.500 ;
        RECT -15.950 22.330 -15.450 22.500 ;
        RECT -15.160 22.330 -14.660 22.500 ;
        RECT -14.370 22.330 -13.870 22.500 ;
        RECT -13.580 22.330 -13.080 22.500 ;
        RECT -12.790 22.330 -12.290 22.500 ;
        RECT -12.000 22.330 -11.500 22.500 ;
        RECT -11.210 22.330 -10.710 22.500 ;
        RECT -10.420 22.330 -9.920 22.500 ;
        RECT -9.630 22.330 -9.130 22.500 ;
        RECT -8.840 22.330 -8.340 22.500 ;
        RECT -8.050 22.330 -7.550 22.500 ;
        RECT -7.260 22.330 -6.760 22.500 ;
        RECT -6.470 22.330 -5.970 22.500 ;
        RECT -5.680 22.330 -5.180 22.500 ;
        RECT -4.890 22.330 -4.390 22.500 ;
        RECT -4.100 22.330 -3.600 22.500 ;
        RECT -3.310 22.330 -2.810 22.500 ;
        RECT -2.520 22.330 -2.020 22.500 ;
        RECT -1.730 22.330 -1.230 22.500 ;
        RECT -0.940 22.330 -0.440 22.500 ;
        RECT -0.150 22.330 0.350 22.500 ;
        RECT 0.640 22.330 1.140 22.500 ;
        RECT 1.430 22.330 1.930 22.500 ;
        RECT 2.220 22.330 2.720 22.500 ;
        RECT 3.010 22.330 3.510 22.500 ;
        RECT 3.800 22.330 4.300 22.500 ;
        RECT 4.590 22.330 5.090 22.500 ;
        RECT 5.380 22.330 5.880 22.500 ;
        RECT 6.170 22.330 6.670 22.500 ;
        RECT 6.960 22.330 7.460 22.500 ;
        RECT 7.750 22.330 8.250 22.500 ;
        RECT 8.540 22.330 9.040 22.500 ;
        RECT 9.330 22.330 9.830 22.500 ;
        RECT 10.120 22.330 10.620 22.500 ;
        RECT 10.910 22.330 11.410 22.500 ;
        RECT -19.900 21.790 -19.400 21.960 ;
        RECT -19.110 21.790 -18.610 21.960 ;
        RECT -18.320 21.790 -17.820 21.960 ;
        RECT -17.530 21.790 -17.030 21.960 ;
        RECT -16.740 21.790 -16.240 21.960 ;
        RECT -15.950 21.790 -15.450 21.960 ;
        RECT -15.160 21.790 -14.660 21.960 ;
        RECT -14.370 21.790 -13.870 21.960 ;
        RECT -13.580 21.790 -13.080 21.960 ;
        RECT -12.790 21.790 -12.290 21.960 ;
        RECT -12.000 21.790 -11.500 21.960 ;
        RECT -11.210 21.790 -10.710 21.960 ;
        RECT -10.420 21.790 -9.920 21.960 ;
        RECT -9.630 21.790 -9.130 21.960 ;
        RECT -8.840 21.790 -8.340 21.960 ;
        RECT -8.050 21.790 -7.550 21.960 ;
        RECT -7.260 21.790 -6.760 21.960 ;
        RECT -6.470 21.790 -5.970 21.960 ;
        RECT -5.680 21.790 -5.180 21.960 ;
        RECT -4.890 21.790 -4.390 21.960 ;
        RECT -4.100 21.790 -3.600 21.960 ;
        RECT -3.310 21.790 -2.810 21.960 ;
        RECT -2.520 21.790 -2.020 21.960 ;
        RECT -1.730 21.790 -1.230 21.960 ;
        RECT -0.940 21.790 -0.440 21.960 ;
        RECT -0.150 21.790 0.350 21.960 ;
        RECT 0.640 21.790 1.140 21.960 ;
        RECT 1.430 21.790 1.930 21.960 ;
        RECT 2.220 21.790 2.720 21.960 ;
        RECT 3.010 21.790 3.510 21.960 ;
        RECT 3.800 21.790 4.300 21.960 ;
        RECT 4.590 21.790 5.090 21.960 ;
        RECT 5.380 21.790 5.880 21.960 ;
        RECT 6.170 21.790 6.670 21.960 ;
        RECT 6.960 21.790 7.460 21.960 ;
        RECT 7.750 21.790 8.250 21.960 ;
        RECT 8.540 21.790 9.040 21.960 ;
        RECT 9.330 21.790 9.830 21.960 ;
        RECT 10.120 21.790 10.620 21.960 ;
        RECT 10.910 21.790 11.410 21.960 ;
        RECT -19.900 20.150 -19.400 20.320 ;
        RECT -19.110 20.150 -18.610 20.320 ;
        RECT -18.320 20.150 -17.820 20.320 ;
        RECT -17.530 20.150 -17.030 20.320 ;
        RECT -16.740 20.150 -16.240 20.320 ;
        RECT -15.950 20.150 -15.450 20.320 ;
        RECT -15.160 20.150 -14.660 20.320 ;
        RECT -14.370 20.150 -13.870 20.320 ;
        RECT -13.580 20.150 -13.080 20.320 ;
        RECT -12.790 20.150 -12.290 20.320 ;
        RECT -12.000 20.150 -11.500 20.320 ;
        RECT -11.210 20.150 -10.710 20.320 ;
        RECT -10.420 20.150 -9.920 20.320 ;
        RECT -9.630 20.150 -9.130 20.320 ;
        RECT -8.840 20.150 -8.340 20.320 ;
        RECT -8.050 20.150 -7.550 20.320 ;
        RECT -7.260 20.150 -6.760 20.320 ;
        RECT -6.470 20.150 -5.970 20.320 ;
        RECT -5.680 20.150 -5.180 20.320 ;
        RECT -4.890 20.150 -4.390 20.320 ;
        RECT -4.100 20.150 -3.600 20.320 ;
        RECT -3.310 20.150 -2.810 20.320 ;
        RECT -2.520 20.150 -2.020 20.320 ;
        RECT -1.730 20.150 -1.230 20.320 ;
        RECT -0.940 20.150 -0.440 20.320 ;
        RECT -0.150 20.150 0.350 20.320 ;
        RECT 0.640 20.150 1.140 20.320 ;
        RECT 1.430 20.150 1.930 20.320 ;
        RECT 2.220 20.150 2.720 20.320 ;
        RECT 3.010 20.150 3.510 20.320 ;
        RECT 3.800 20.150 4.300 20.320 ;
        RECT 4.590 20.150 5.090 20.320 ;
        RECT 5.380 20.150 5.880 20.320 ;
        RECT 6.170 20.150 6.670 20.320 ;
        RECT 6.960 20.150 7.460 20.320 ;
        RECT 7.750 20.150 8.250 20.320 ;
        RECT 8.540 20.150 9.040 20.320 ;
        RECT 9.330 20.150 9.830 20.320 ;
        RECT 10.120 20.150 10.620 20.320 ;
        RECT 10.910 20.150 11.410 20.320 ;
        RECT -19.900 18.770 -19.400 18.940 ;
        RECT -19.110 18.770 -18.610 18.940 ;
        RECT -18.320 18.770 -17.820 18.940 ;
        RECT -17.530 18.770 -17.030 18.940 ;
        RECT -16.740 18.770 -16.240 18.940 ;
        RECT -15.950 18.770 -15.450 18.940 ;
        RECT -15.160 18.770 -14.660 18.940 ;
        RECT -14.370 18.770 -13.870 18.940 ;
        RECT -13.580 18.770 -13.080 18.940 ;
        RECT -12.790 18.770 -12.290 18.940 ;
        RECT -12.000 18.770 -11.500 18.940 ;
        RECT -11.210 18.770 -10.710 18.940 ;
        RECT -10.420 18.770 -9.920 18.940 ;
        RECT -9.630 18.770 -9.130 18.940 ;
        RECT -8.840 18.770 -8.340 18.940 ;
        RECT -8.050 18.770 -7.550 18.940 ;
        RECT -7.260 18.770 -6.760 18.940 ;
        RECT -6.470 18.770 -5.970 18.940 ;
        RECT -5.680 18.770 -5.180 18.940 ;
        RECT -4.890 18.770 -4.390 18.940 ;
        RECT -4.100 18.770 -3.600 18.940 ;
        RECT -3.310 18.770 -2.810 18.940 ;
        RECT -2.520 18.770 -2.020 18.940 ;
        RECT -1.730 18.770 -1.230 18.940 ;
        RECT -0.940 18.770 -0.440 18.940 ;
        RECT -0.150 18.770 0.350 18.940 ;
        RECT 0.640 18.770 1.140 18.940 ;
        RECT 1.430 18.770 1.930 18.940 ;
        RECT 2.220 18.770 2.720 18.940 ;
        RECT 3.010 18.770 3.510 18.940 ;
        RECT 3.800 18.770 4.300 18.940 ;
        RECT 4.590 18.770 5.090 18.940 ;
        RECT 5.380 18.770 5.880 18.940 ;
        RECT 6.170 18.770 6.670 18.940 ;
        RECT 6.960 18.770 7.460 18.940 ;
        RECT 7.750 18.770 8.250 18.940 ;
        RECT 8.540 18.770 9.040 18.940 ;
        RECT 9.330 18.770 9.830 18.940 ;
        RECT 10.120 18.770 10.620 18.940 ;
        RECT 10.910 18.770 11.410 18.940 ;
        RECT -19.900 17.130 -19.400 17.300 ;
        RECT -19.110 17.130 -18.610 17.300 ;
        RECT -18.320 17.130 -17.820 17.300 ;
        RECT -17.530 17.130 -17.030 17.300 ;
        RECT -16.740 17.130 -16.240 17.300 ;
        RECT -15.950 17.130 -15.450 17.300 ;
        RECT -15.160 17.130 -14.660 17.300 ;
        RECT -14.370 17.130 -13.870 17.300 ;
        RECT -13.580 17.130 -13.080 17.300 ;
        RECT -12.790 17.130 -12.290 17.300 ;
        RECT -12.000 17.130 -11.500 17.300 ;
        RECT -11.210 17.130 -10.710 17.300 ;
        RECT -10.420 17.130 -9.920 17.300 ;
        RECT -9.630 17.130 -9.130 17.300 ;
        RECT -8.840 17.130 -8.340 17.300 ;
        RECT -8.050 17.130 -7.550 17.300 ;
        RECT -7.260 17.130 -6.760 17.300 ;
        RECT -6.470 17.130 -5.970 17.300 ;
        RECT -5.680 17.130 -5.180 17.300 ;
        RECT -4.890 17.130 -4.390 17.300 ;
        RECT -4.100 17.130 -3.600 17.300 ;
        RECT -3.310 17.130 -2.810 17.300 ;
        RECT -2.520 17.130 -2.020 17.300 ;
        RECT -1.730 17.130 -1.230 17.300 ;
        RECT -0.940 17.130 -0.440 17.300 ;
        RECT -0.150 17.130 0.350 17.300 ;
        RECT 0.640 17.130 1.140 17.300 ;
        RECT 1.430 17.130 1.930 17.300 ;
        RECT 2.220 17.130 2.720 17.300 ;
        RECT 3.010 17.130 3.510 17.300 ;
        RECT 3.800 17.130 4.300 17.300 ;
        RECT 4.590 17.130 5.090 17.300 ;
        RECT 5.380 17.130 5.880 17.300 ;
        RECT 6.170 17.130 6.670 17.300 ;
        RECT 6.960 17.130 7.460 17.300 ;
        RECT 7.750 17.130 8.250 17.300 ;
        RECT 8.540 17.130 9.040 17.300 ;
        RECT 9.330 17.130 9.830 17.300 ;
        RECT 10.120 17.130 10.620 17.300 ;
        RECT 10.910 17.130 11.410 17.300 ;
        RECT -19.900 16.590 -19.400 16.760 ;
        RECT -19.110 16.590 -18.610 16.760 ;
        RECT -18.320 16.590 -17.820 16.760 ;
        RECT -17.530 16.590 -17.030 16.760 ;
        RECT -16.740 16.590 -16.240 16.760 ;
        RECT -15.950 16.590 -15.450 16.760 ;
        RECT -15.160 16.590 -14.660 16.760 ;
        RECT -14.370 16.590 -13.870 16.760 ;
        RECT -13.580 16.590 -13.080 16.760 ;
        RECT -12.790 16.590 -12.290 16.760 ;
        RECT -12.000 16.590 -11.500 16.760 ;
        RECT -11.210 16.590 -10.710 16.760 ;
        RECT -10.420 16.590 -9.920 16.760 ;
        RECT -9.630 16.590 -9.130 16.760 ;
        RECT -8.840 16.590 -8.340 16.760 ;
        RECT -8.050 16.590 -7.550 16.760 ;
        RECT -7.260 16.590 -6.760 16.760 ;
        RECT -6.470 16.590 -5.970 16.760 ;
        RECT -5.680 16.590 -5.180 16.760 ;
        RECT -4.890 16.590 -4.390 16.760 ;
        RECT -4.100 16.590 -3.600 16.760 ;
        RECT -3.310 16.590 -2.810 16.760 ;
        RECT -2.520 16.590 -2.020 16.760 ;
        RECT -1.730 16.590 -1.230 16.760 ;
        RECT -0.940 16.590 -0.440 16.760 ;
        RECT -0.150 16.590 0.350 16.760 ;
        RECT 0.640 16.590 1.140 16.760 ;
        RECT 1.430 16.590 1.930 16.760 ;
        RECT 2.220 16.590 2.720 16.760 ;
        RECT 3.010 16.590 3.510 16.760 ;
        RECT 3.800 16.590 4.300 16.760 ;
        RECT 4.590 16.590 5.090 16.760 ;
        RECT 5.380 16.590 5.880 16.760 ;
        RECT 6.170 16.590 6.670 16.760 ;
        RECT 6.960 16.590 7.460 16.760 ;
        RECT 7.750 16.590 8.250 16.760 ;
        RECT 8.540 16.590 9.040 16.760 ;
        RECT 9.330 16.590 9.830 16.760 ;
        RECT 10.120 16.590 10.620 16.760 ;
        RECT 10.910 16.590 11.410 16.760 ;
        RECT -19.900 14.950 -19.400 15.120 ;
        RECT -19.110 14.950 -18.610 15.120 ;
        RECT -18.320 14.950 -17.820 15.120 ;
        RECT -17.530 14.950 -17.030 15.120 ;
        RECT -16.740 14.950 -16.240 15.120 ;
        RECT -15.950 14.950 -15.450 15.120 ;
        RECT -15.160 14.950 -14.660 15.120 ;
        RECT -14.370 14.950 -13.870 15.120 ;
        RECT -13.580 14.950 -13.080 15.120 ;
        RECT -12.790 14.950 -12.290 15.120 ;
        RECT -12.000 14.950 -11.500 15.120 ;
        RECT -11.210 14.950 -10.710 15.120 ;
        RECT -10.420 14.950 -9.920 15.120 ;
        RECT -9.630 14.950 -9.130 15.120 ;
        RECT -8.840 14.950 -8.340 15.120 ;
        RECT -8.050 14.950 -7.550 15.120 ;
        RECT -7.260 14.950 -6.760 15.120 ;
        RECT -6.470 14.950 -5.970 15.120 ;
        RECT -5.680 14.950 -5.180 15.120 ;
        RECT -4.890 14.950 -4.390 15.120 ;
        RECT -4.100 14.950 -3.600 15.120 ;
        RECT -3.310 14.950 -2.810 15.120 ;
        RECT -2.520 14.950 -2.020 15.120 ;
        RECT -1.730 14.950 -1.230 15.120 ;
        RECT -0.940 14.950 -0.440 15.120 ;
        RECT -0.150 14.950 0.350 15.120 ;
        RECT 0.640 14.950 1.140 15.120 ;
        RECT 1.430 14.950 1.930 15.120 ;
        RECT 2.220 14.950 2.720 15.120 ;
        RECT 3.010 14.950 3.510 15.120 ;
        RECT 3.800 14.950 4.300 15.120 ;
        RECT 4.590 14.950 5.090 15.120 ;
        RECT 5.380 14.950 5.880 15.120 ;
        RECT 6.170 14.950 6.670 15.120 ;
        RECT 6.960 14.950 7.460 15.120 ;
        RECT 7.750 14.950 8.250 15.120 ;
        RECT 8.540 14.950 9.040 15.120 ;
        RECT 9.330 14.950 9.830 15.120 ;
        RECT 10.120 14.950 10.620 15.120 ;
        RECT 10.910 14.950 11.410 15.120 ;
        RECT -19.900 14.410 -19.400 14.580 ;
        RECT -19.110 14.410 -18.610 14.580 ;
        RECT -18.320 14.410 -17.820 14.580 ;
        RECT -17.530 14.410 -17.030 14.580 ;
        RECT -16.740 14.410 -16.240 14.580 ;
        RECT -15.950 14.410 -15.450 14.580 ;
        RECT -15.160 14.410 -14.660 14.580 ;
        RECT -14.370 14.410 -13.870 14.580 ;
        RECT -13.580 14.410 -13.080 14.580 ;
        RECT -12.790 14.410 -12.290 14.580 ;
        RECT -12.000 14.410 -11.500 14.580 ;
        RECT -11.210 14.410 -10.710 14.580 ;
        RECT -10.420 14.410 -9.920 14.580 ;
        RECT -9.630 14.410 -9.130 14.580 ;
        RECT -8.840 14.410 -8.340 14.580 ;
        RECT -8.050 14.410 -7.550 14.580 ;
        RECT -7.260 14.410 -6.760 14.580 ;
        RECT -6.470 14.410 -5.970 14.580 ;
        RECT -5.680 14.410 -5.180 14.580 ;
        RECT -4.890 14.410 -4.390 14.580 ;
        RECT -4.100 14.410 -3.600 14.580 ;
        RECT -3.310 14.410 -2.810 14.580 ;
        RECT -2.520 14.410 -2.020 14.580 ;
        RECT -1.730 14.410 -1.230 14.580 ;
        RECT -0.940 14.410 -0.440 14.580 ;
        RECT -0.150 14.410 0.350 14.580 ;
        RECT 0.640 14.410 1.140 14.580 ;
        RECT 1.430 14.410 1.930 14.580 ;
        RECT 2.220 14.410 2.720 14.580 ;
        RECT 3.010 14.410 3.510 14.580 ;
        RECT 3.800 14.410 4.300 14.580 ;
        RECT 4.590 14.410 5.090 14.580 ;
        RECT 5.380 14.410 5.880 14.580 ;
        RECT 6.170 14.410 6.670 14.580 ;
        RECT 6.960 14.410 7.460 14.580 ;
        RECT 7.750 14.410 8.250 14.580 ;
        RECT 8.540 14.410 9.040 14.580 ;
        RECT 9.330 14.410 9.830 14.580 ;
        RECT 10.120 14.410 10.620 14.580 ;
        RECT 10.910 14.410 11.410 14.580 ;
        RECT -19.900 12.770 -19.400 12.940 ;
        RECT -19.110 12.770 -18.610 12.940 ;
        RECT -18.320 12.770 -17.820 12.940 ;
        RECT -17.530 12.770 -17.030 12.940 ;
        RECT -16.740 12.770 -16.240 12.940 ;
        RECT -15.950 12.770 -15.450 12.940 ;
        RECT -15.160 12.770 -14.660 12.940 ;
        RECT -14.370 12.770 -13.870 12.940 ;
        RECT -13.580 12.770 -13.080 12.940 ;
        RECT -12.790 12.770 -12.290 12.940 ;
        RECT -12.000 12.770 -11.500 12.940 ;
        RECT -11.210 12.770 -10.710 12.940 ;
        RECT -10.420 12.770 -9.920 12.940 ;
        RECT -9.630 12.770 -9.130 12.940 ;
        RECT -8.840 12.770 -8.340 12.940 ;
        RECT -8.050 12.770 -7.550 12.940 ;
        RECT -7.260 12.770 -6.760 12.940 ;
        RECT -6.470 12.770 -5.970 12.940 ;
        RECT -5.680 12.770 -5.180 12.940 ;
        RECT -4.890 12.770 -4.390 12.940 ;
        RECT -4.100 12.770 -3.600 12.940 ;
        RECT -3.310 12.770 -2.810 12.940 ;
        RECT -2.520 12.770 -2.020 12.940 ;
        RECT -1.730 12.770 -1.230 12.940 ;
        RECT -0.940 12.770 -0.440 12.940 ;
        RECT -0.150 12.770 0.350 12.940 ;
        RECT 0.640 12.770 1.140 12.940 ;
        RECT 1.430 12.770 1.930 12.940 ;
        RECT 2.220 12.770 2.720 12.940 ;
        RECT 3.010 12.770 3.510 12.940 ;
        RECT 3.800 12.770 4.300 12.940 ;
        RECT 4.590 12.770 5.090 12.940 ;
        RECT 5.380 12.770 5.880 12.940 ;
        RECT 6.170 12.770 6.670 12.940 ;
        RECT 6.960 12.770 7.460 12.940 ;
        RECT 7.750 12.770 8.250 12.940 ;
        RECT 8.540 12.770 9.040 12.940 ;
        RECT 9.330 12.770 9.830 12.940 ;
        RECT 10.120 12.770 10.620 12.940 ;
        RECT 10.910 12.770 11.410 12.940 ;
        RECT -19.900 12.230 -19.400 12.400 ;
        RECT -19.110 12.230 -18.610 12.400 ;
        RECT -18.320 12.230 -17.820 12.400 ;
        RECT -17.530 12.230 -17.030 12.400 ;
        RECT -16.740 12.230 -16.240 12.400 ;
        RECT -15.950 12.230 -15.450 12.400 ;
        RECT -15.160 12.230 -14.660 12.400 ;
        RECT -14.370 12.230 -13.870 12.400 ;
        RECT -13.580 12.230 -13.080 12.400 ;
        RECT -12.790 12.230 -12.290 12.400 ;
        RECT -12.000 12.230 -11.500 12.400 ;
        RECT -11.210 12.230 -10.710 12.400 ;
        RECT -10.420 12.230 -9.920 12.400 ;
        RECT -9.630 12.230 -9.130 12.400 ;
        RECT -8.840 12.230 -8.340 12.400 ;
        RECT -8.050 12.230 -7.550 12.400 ;
        RECT -7.260 12.230 -6.760 12.400 ;
        RECT -6.470 12.230 -5.970 12.400 ;
        RECT -5.680 12.230 -5.180 12.400 ;
        RECT -4.890 12.230 -4.390 12.400 ;
        RECT -4.100 12.230 -3.600 12.400 ;
        RECT -3.310 12.230 -2.810 12.400 ;
        RECT -2.520 12.230 -2.020 12.400 ;
        RECT -1.730 12.230 -1.230 12.400 ;
        RECT -0.940 12.230 -0.440 12.400 ;
        RECT -0.150 12.230 0.350 12.400 ;
        RECT 0.640 12.230 1.140 12.400 ;
        RECT 1.430 12.230 1.930 12.400 ;
        RECT 2.220 12.230 2.720 12.400 ;
        RECT 3.010 12.230 3.510 12.400 ;
        RECT 3.800 12.230 4.300 12.400 ;
        RECT 4.590 12.230 5.090 12.400 ;
        RECT 5.380 12.230 5.880 12.400 ;
        RECT 6.170 12.230 6.670 12.400 ;
        RECT 6.960 12.230 7.460 12.400 ;
        RECT 7.750 12.230 8.250 12.400 ;
        RECT 8.540 12.230 9.040 12.400 ;
        RECT 9.330 12.230 9.830 12.400 ;
        RECT 10.120 12.230 10.620 12.400 ;
        RECT 10.910 12.230 11.410 12.400 ;
        RECT -19.900 10.590 -19.400 10.760 ;
        RECT -19.110 10.590 -18.610 10.760 ;
        RECT -18.320 10.590 -17.820 10.760 ;
        RECT -17.530 10.590 -17.030 10.760 ;
        RECT -16.740 10.590 -16.240 10.760 ;
        RECT -15.950 10.590 -15.450 10.760 ;
        RECT -15.160 10.590 -14.660 10.760 ;
        RECT -14.370 10.590 -13.870 10.760 ;
        RECT -13.580 10.590 -13.080 10.760 ;
        RECT -12.790 10.590 -12.290 10.760 ;
        RECT -12.000 10.590 -11.500 10.760 ;
        RECT -11.210 10.590 -10.710 10.760 ;
        RECT -10.420 10.590 -9.920 10.760 ;
        RECT -9.630 10.590 -9.130 10.760 ;
        RECT -8.840 10.590 -8.340 10.760 ;
        RECT -8.050 10.590 -7.550 10.760 ;
        RECT -7.260 10.590 -6.760 10.760 ;
        RECT -6.470 10.590 -5.970 10.760 ;
        RECT -5.680 10.590 -5.180 10.760 ;
        RECT -4.890 10.590 -4.390 10.760 ;
        RECT -4.100 10.590 -3.600 10.760 ;
        RECT -3.310 10.590 -2.810 10.760 ;
        RECT -2.520 10.590 -2.020 10.760 ;
        RECT -1.730 10.590 -1.230 10.760 ;
        RECT -0.940 10.590 -0.440 10.760 ;
        RECT -0.150 10.590 0.350 10.760 ;
        RECT 0.640 10.590 1.140 10.760 ;
        RECT 1.430 10.590 1.930 10.760 ;
        RECT 2.220 10.590 2.720 10.760 ;
        RECT 3.010 10.590 3.510 10.760 ;
        RECT 3.800 10.590 4.300 10.760 ;
        RECT 4.590 10.590 5.090 10.760 ;
        RECT 5.380 10.590 5.880 10.760 ;
        RECT 6.170 10.590 6.670 10.760 ;
        RECT 6.960 10.590 7.460 10.760 ;
        RECT 7.750 10.590 8.250 10.760 ;
        RECT 8.540 10.590 9.040 10.760 ;
        RECT 9.330 10.590 9.830 10.760 ;
        RECT 10.120 10.590 10.620 10.760 ;
        RECT 10.910 10.590 11.410 10.760 ;
        RECT -19.900 10.050 -19.400 10.220 ;
        RECT -19.110 10.050 -18.610 10.220 ;
        RECT -18.320 10.050 -17.820 10.220 ;
        RECT -17.530 10.050 -17.030 10.220 ;
        RECT -16.740 10.050 -16.240 10.220 ;
        RECT -15.950 10.050 -15.450 10.220 ;
        RECT -15.160 10.050 -14.660 10.220 ;
        RECT -14.370 10.050 -13.870 10.220 ;
        RECT -13.580 10.050 -13.080 10.220 ;
        RECT -12.790 10.050 -12.290 10.220 ;
        RECT -12.000 10.050 -11.500 10.220 ;
        RECT -11.210 10.050 -10.710 10.220 ;
        RECT -10.420 10.050 -9.920 10.220 ;
        RECT -9.630 10.050 -9.130 10.220 ;
        RECT -8.840 10.050 -8.340 10.220 ;
        RECT -8.050 10.050 -7.550 10.220 ;
        RECT -7.260 10.050 -6.760 10.220 ;
        RECT -6.470 10.050 -5.970 10.220 ;
        RECT -5.680 10.050 -5.180 10.220 ;
        RECT -4.890 10.050 -4.390 10.220 ;
        RECT -4.100 10.050 -3.600 10.220 ;
        RECT -3.310 10.050 -2.810 10.220 ;
        RECT -2.520 10.050 -2.020 10.220 ;
        RECT -1.730 10.050 -1.230 10.220 ;
        RECT -0.940 10.050 -0.440 10.220 ;
        RECT -0.150 10.050 0.350 10.220 ;
        RECT 0.640 10.050 1.140 10.220 ;
        RECT 1.430 10.050 1.930 10.220 ;
        RECT 2.220 10.050 2.720 10.220 ;
        RECT 3.010 10.050 3.510 10.220 ;
        RECT 3.800 10.050 4.300 10.220 ;
        RECT 4.590 10.050 5.090 10.220 ;
        RECT 5.380 10.050 5.880 10.220 ;
        RECT 6.170 10.050 6.670 10.220 ;
        RECT 6.960 10.050 7.460 10.220 ;
        RECT 7.750 10.050 8.250 10.220 ;
        RECT 8.540 10.050 9.040 10.220 ;
        RECT 9.330 10.050 9.830 10.220 ;
        RECT 10.120 10.050 10.620 10.220 ;
        RECT 10.910 10.050 11.410 10.220 ;
        RECT -19.900 8.410 -19.400 8.580 ;
        RECT -19.110 8.410 -18.610 8.580 ;
        RECT -18.320 8.410 -17.820 8.580 ;
        RECT -17.530 8.410 -17.030 8.580 ;
        RECT -16.740 8.410 -16.240 8.580 ;
        RECT -15.950 8.410 -15.450 8.580 ;
        RECT -15.160 8.410 -14.660 8.580 ;
        RECT -14.370 8.410 -13.870 8.580 ;
        RECT -13.580 8.410 -13.080 8.580 ;
        RECT -12.790 8.410 -12.290 8.580 ;
        RECT -12.000 8.410 -11.500 8.580 ;
        RECT -11.210 8.410 -10.710 8.580 ;
        RECT -10.420 8.410 -9.920 8.580 ;
        RECT -9.630 8.410 -9.130 8.580 ;
        RECT -8.840 8.410 -8.340 8.580 ;
        RECT -8.050 8.410 -7.550 8.580 ;
        RECT -7.260 8.410 -6.760 8.580 ;
        RECT -6.470 8.410 -5.970 8.580 ;
        RECT -5.680 8.410 -5.180 8.580 ;
        RECT -4.890 8.410 -4.390 8.580 ;
        RECT -4.100 8.410 -3.600 8.580 ;
        RECT -3.310 8.410 -2.810 8.580 ;
        RECT -2.520 8.410 -2.020 8.580 ;
        RECT -1.730 8.410 -1.230 8.580 ;
        RECT -0.940 8.410 -0.440 8.580 ;
        RECT -0.150 8.410 0.350 8.580 ;
        RECT 0.640 8.410 1.140 8.580 ;
        RECT 1.430 8.410 1.930 8.580 ;
        RECT 2.220 8.410 2.720 8.580 ;
        RECT 3.010 8.410 3.510 8.580 ;
        RECT 3.800 8.410 4.300 8.580 ;
        RECT 4.590 8.410 5.090 8.580 ;
        RECT 5.380 8.410 5.880 8.580 ;
        RECT 6.170 8.410 6.670 8.580 ;
        RECT 6.960 8.410 7.460 8.580 ;
        RECT 7.750 8.410 8.250 8.580 ;
        RECT 8.540 8.410 9.040 8.580 ;
        RECT 9.330 8.410 9.830 8.580 ;
        RECT 10.120 8.410 10.620 8.580 ;
        RECT 10.910 8.410 11.410 8.580 ;
        RECT -15.390 3.180 -15.220 4.220 ;
        RECT -13.810 3.180 -13.640 4.220 ;
        RECT -12.470 3.180 -12.300 4.220 ;
        RECT -10.890 3.180 -10.720 4.220 ;
        RECT -9.550 3.180 -9.380 4.220 ;
        RECT -7.970 3.180 -7.800 4.220 ;
        RECT -6.630 3.180 -6.460 4.220 ;
        RECT -5.050 3.180 -4.880 4.220 ;
        RECT -3.710 3.180 -3.540 4.220 ;
        RECT -2.920 3.180 -2.750 4.220 ;
        RECT -2.130 3.180 -1.960 4.220 ;
        RECT -0.790 3.180 -0.620 4.220 ;
        RECT 0.000 3.180 0.170 4.220 ;
        RECT 0.790 3.180 0.960 4.220 ;
        RECT 2.130 3.180 2.300 4.220 ;
        RECT 3.710 3.180 3.880 4.220 ;
        RECT 5.840 3.180 6.010 4.220 ;
        RECT -15.160 2.795 -14.660 2.965 ;
        RECT -14.370 2.795 -13.870 2.965 ;
        RECT -12.240 2.795 -11.740 2.965 ;
        RECT -11.450 2.795 -10.950 2.965 ;
        RECT -9.320 2.795 -8.820 2.965 ;
        RECT -8.530 2.795 -8.030 2.965 ;
        RECT -6.400 2.795 -5.900 2.965 ;
        RECT -5.610 2.795 -5.110 2.965 ;
        RECT 2.360 2.795 2.860 2.965 ;
        RECT 3.150 2.795 3.650 2.965 ;
        RECT 5.280 2.795 5.780 2.965 ;
        RECT -11.435 -0.095 -10.935 0.075 ;
        RECT -4.925 -0.095 -4.425 0.075 ;
        RECT -2.755 -0.095 -2.255 0.075 ;
        RECT -0.585 -0.095 -0.085 0.075 ;
        RECT 1.580 -0.100 2.080 0.070 ;
        RECT 2.370 -0.100 2.870 0.070 ;
        RECT 3.160 -0.100 3.660 0.070 ;
        RECT 3.950 -0.100 4.450 0.070 ;
        RECT 6.125 -0.095 6.625 0.075 ;
        RECT -16.005 -1.305 -15.835 -0.265 ;
        RECT -15.215 -1.305 -15.045 -0.265 ;
        RECT -13.835 -1.305 -13.665 -0.265 ;
        RECT -13.045 -1.305 -12.875 -0.265 ;
        RECT -10.875 -1.305 -10.705 -0.265 ;
        RECT -9.495 -1.305 -9.325 -0.265 ;
        RECT -8.705 -1.305 -8.535 -0.265 ;
        RECT -7.325 -1.305 -7.155 -0.265 ;
        RECT -6.535 -1.305 -6.365 -0.265 ;
        RECT -4.365 -1.305 -4.195 -0.265 ;
        RECT -2.985 -1.305 -2.815 -0.265 ;
        RECT -0.025 -1.305 0.145 -0.265 ;
        RECT 2.140 -1.310 2.310 -0.270 ;
        RECT 3.720 -1.310 3.890 -0.270 ;
        RECT 5.895 -1.305 6.065 -0.265 ;
        RECT 8.070 -1.305 8.240 -0.265 ;
        RECT 8.860 -1.305 9.030 -0.265 ;
        RECT -11.435 -1.645 -10.935 -1.475 ;
        RECT -4.925 -1.645 -4.425 -1.475 ;
        RECT -2.755 -1.645 -2.255 -1.475 ;
        RECT -0.585 -1.645 -0.085 -1.475 ;
        RECT 1.580 -1.650 2.080 -1.480 ;
        RECT 2.370 -1.650 2.870 -1.480 ;
        RECT 3.160 -1.650 3.660 -1.480 ;
        RECT 3.950 -1.650 4.450 -1.480 ;
        RECT 6.125 -1.645 6.625 -1.475 ;
        RECT -19.980 -4.180 -19.480 -4.010 ;
        RECT -19.190 -4.180 -18.690 -4.010 ;
        RECT -18.400 -4.180 -17.900 -4.010 ;
        RECT -17.610 -4.180 -17.110 -4.010 ;
        RECT -16.820 -4.180 -16.320 -4.010 ;
        RECT -16.030 -4.180 -15.530 -4.010 ;
        RECT -15.240 -4.180 -14.740 -4.010 ;
        RECT -14.450 -4.180 -13.950 -4.010 ;
        RECT -13.660 -4.180 -13.160 -4.010 ;
        RECT -12.870 -4.180 -12.370 -4.010 ;
        RECT -12.080 -4.180 -11.580 -4.010 ;
        RECT -11.290 -4.180 -10.790 -4.010 ;
        RECT -10.500 -4.180 -10.000 -4.010 ;
        RECT -9.710 -4.180 -9.210 -4.010 ;
        RECT -8.920 -4.180 -8.420 -4.010 ;
        RECT -8.130 -4.180 -7.630 -4.010 ;
        RECT -7.340 -4.180 -6.840 -4.010 ;
        RECT -6.550 -4.180 -6.050 -4.010 ;
        RECT -5.760 -4.180 -5.260 -4.010 ;
        RECT -4.970 -4.180 -4.470 -4.010 ;
        RECT -4.180 -4.180 -3.680 -4.010 ;
        RECT -3.390 -4.180 -2.890 -4.010 ;
        RECT -2.600 -4.180 -2.100 -4.010 ;
        RECT -1.810 -4.180 -1.310 -4.010 ;
        RECT -1.020 -4.180 -0.520 -4.010 ;
        RECT -0.230 -4.180 0.270 -4.010 ;
        RECT 0.560 -4.180 1.060 -4.010 ;
        RECT 1.350 -4.180 1.850 -4.010 ;
        RECT 2.140 -4.180 2.640 -4.010 ;
        RECT 2.930 -4.180 3.430 -4.010 ;
        RECT 3.720 -4.180 4.220 -4.010 ;
        RECT 4.510 -4.180 5.010 -4.010 ;
        RECT 5.300 -4.180 5.800 -4.010 ;
        RECT 6.090 -4.180 6.590 -4.010 ;
        RECT 6.880 -4.180 7.380 -4.010 ;
        RECT 7.670 -4.180 8.170 -4.010 ;
        RECT 8.460 -4.180 8.960 -4.010 ;
        RECT 9.250 -4.180 9.750 -4.010 ;
        RECT 10.040 -4.180 10.540 -4.010 ;
        RECT 10.830 -4.180 11.330 -4.010 ;
        RECT -19.980 -5.730 -19.480 -5.560 ;
        RECT -19.190 -5.730 -18.690 -5.560 ;
        RECT -18.400 -5.730 -17.900 -5.560 ;
        RECT -17.610 -5.730 -17.110 -5.560 ;
        RECT -16.820 -5.730 -16.320 -5.560 ;
        RECT -16.030 -5.730 -15.530 -5.560 ;
        RECT -15.240 -5.730 -14.740 -5.560 ;
        RECT -14.450 -5.730 -13.950 -5.560 ;
        RECT -13.660 -5.730 -13.160 -5.560 ;
        RECT -12.870 -5.730 -12.370 -5.560 ;
        RECT -12.080 -5.730 -11.580 -5.560 ;
        RECT -11.290 -5.730 -10.790 -5.560 ;
        RECT -10.500 -5.730 -10.000 -5.560 ;
        RECT -9.710 -5.730 -9.210 -5.560 ;
        RECT -8.920 -5.730 -8.420 -5.560 ;
        RECT -8.130 -5.730 -7.630 -5.560 ;
        RECT -7.340 -5.730 -6.840 -5.560 ;
        RECT -6.550 -5.730 -6.050 -5.560 ;
        RECT -5.760 -5.730 -5.260 -5.560 ;
        RECT -4.970 -5.730 -4.470 -5.560 ;
        RECT -4.180 -5.730 -3.680 -5.560 ;
        RECT -3.390 -5.730 -2.890 -5.560 ;
        RECT -2.600 -5.730 -2.100 -5.560 ;
        RECT -1.810 -5.730 -1.310 -5.560 ;
        RECT -1.020 -5.730 -0.520 -5.560 ;
        RECT -0.230 -5.730 0.270 -5.560 ;
        RECT 0.560 -5.730 1.060 -5.560 ;
        RECT 1.350 -5.730 1.850 -5.560 ;
        RECT 2.140 -5.730 2.640 -5.560 ;
        RECT 2.930 -5.730 3.430 -5.560 ;
        RECT 3.720 -5.730 4.220 -5.560 ;
        RECT 4.510 -5.730 5.010 -5.560 ;
        RECT 5.300 -5.730 5.800 -5.560 ;
        RECT 6.090 -5.730 6.590 -5.560 ;
        RECT 6.880 -5.730 7.380 -5.560 ;
        RECT 7.670 -5.730 8.170 -5.560 ;
        RECT 8.460 -5.730 8.960 -5.560 ;
        RECT 9.250 -5.730 9.750 -5.560 ;
        RECT 10.040 -5.730 10.540 -5.560 ;
        RECT 10.830 -5.730 11.330 -5.560 ;
        RECT -19.980 -6.270 -19.480 -6.100 ;
        RECT -19.190 -6.270 -18.690 -6.100 ;
        RECT -18.400 -6.270 -17.900 -6.100 ;
        RECT -17.610 -6.270 -17.110 -6.100 ;
        RECT -16.820 -6.270 -16.320 -6.100 ;
        RECT -16.030 -6.270 -15.530 -6.100 ;
        RECT -15.240 -6.270 -14.740 -6.100 ;
        RECT -14.450 -6.270 -13.950 -6.100 ;
        RECT -13.660 -6.270 -13.160 -6.100 ;
        RECT -12.870 -6.270 -12.370 -6.100 ;
        RECT -12.080 -6.270 -11.580 -6.100 ;
        RECT -11.290 -6.270 -10.790 -6.100 ;
        RECT -10.500 -6.270 -10.000 -6.100 ;
        RECT -9.710 -6.270 -9.210 -6.100 ;
        RECT -8.920 -6.270 -8.420 -6.100 ;
        RECT -8.130 -6.270 -7.630 -6.100 ;
        RECT -7.340 -6.270 -6.840 -6.100 ;
        RECT -6.550 -6.270 -6.050 -6.100 ;
        RECT -5.760 -6.270 -5.260 -6.100 ;
        RECT -4.970 -6.270 -4.470 -6.100 ;
        RECT -4.180 -6.270 -3.680 -6.100 ;
        RECT -3.390 -6.270 -2.890 -6.100 ;
        RECT -2.600 -6.270 -2.100 -6.100 ;
        RECT -1.810 -6.270 -1.310 -6.100 ;
        RECT -1.020 -6.270 -0.520 -6.100 ;
        RECT -0.230 -6.270 0.270 -6.100 ;
        RECT 0.560 -6.270 1.060 -6.100 ;
        RECT 1.350 -6.270 1.850 -6.100 ;
        RECT 2.140 -6.270 2.640 -6.100 ;
        RECT 2.930 -6.270 3.430 -6.100 ;
        RECT 3.720 -6.270 4.220 -6.100 ;
        RECT 4.510 -6.270 5.010 -6.100 ;
        RECT 5.300 -6.270 5.800 -6.100 ;
        RECT 6.090 -6.270 6.590 -6.100 ;
        RECT 6.880 -6.270 7.380 -6.100 ;
        RECT 7.670 -6.270 8.170 -6.100 ;
        RECT 8.460 -6.270 8.960 -6.100 ;
        RECT 9.250 -6.270 9.750 -6.100 ;
        RECT 10.040 -6.270 10.540 -6.100 ;
        RECT 10.830 -6.270 11.330 -6.100 ;
        RECT -19.980 -7.820 -19.480 -7.650 ;
        RECT -19.190 -7.820 -18.690 -7.650 ;
        RECT -18.400 -7.820 -17.900 -7.650 ;
        RECT -17.610 -7.820 -17.110 -7.650 ;
        RECT -16.820 -7.820 -16.320 -7.650 ;
        RECT -16.030 -7.820 -15.530 -7.650 ;
        RECT -15.240 -7.820 -14.740 -7.650 ;
        RECT -14.450 -7.820 -13.950 -7.650 ;
        RECT -13.660 -7.820 -13.160 -7.650 ;
        RECT -12.870 -7.820 -12.370 -7.650 ;
        RECT -12.080 -7.820 -11.580 -7.650 ;
        RECT -11.290 -7.820 -10.790 -7.650 ;
        RECT -10.500 -7.820 -10.000 -7.650 ;
        RECT -9.710 -7.820 -9.210 -7.650 ;
        RECT -8.920 -7.820 -8.420 -7.650 ;
        RECT -8.130 -7.820 -7.630 -7.650 ;
        RECT -7.340 -7.820 -6.840 -7.650 ;
        RECT -6.550 -7.820 -6.050 -7.650 ;
        RECT -5.760 -7.820 -5.260 -7.650 ;
        RECT -4.970 -7.820 -4.470 -7.650 ;
        RECT -4.180 -7.820 -3.680 -7.650 ;
        RECT -3.390 -7.820 -2.890 -7.650 ;
        RECT -2.600 -7.820 -2.100 -7.650 ;
        RECT -1.810 -7.820 -1.310 -7.650 ;
        RECT -1.020 -7.820 -0.520 -7.650 ;
        RECT -0.230 -7.820 0.270 -7.650 ;
        RECT 0.560 -7.820 1.060 -7.650 ;
        RECT 1.350 -7.820 1.850 -7.650 ;
        RECT 2.140 -7.820 2.640 -7.650 ;
        RECT 2.930 -7.820 3.430 -7.650 ;
        RECT 3.720 -7.820 4.220 -7.650 ;
        RECT 4.510 -7.820 5.010 -7.650 ;
        RECT 5.300 -7.820 5.800 -7.650 ;
        RECT 6.090 -7.820 6.590 -7.650 ;
        RECT 6.880 -7.820 7.380 -7.650 ;
        RECT 7.670 -7.820 8.170 -7.650 ;
        RECT 8.460 -7.820 8.960 -7.650 ;
        RECT 9.250 -7.820 9.750 -7.650 ;
        RECT 10.040 -7.820 10.540 -7.650 ;
        RECT 10.830 -7.820 11.330 -7.650 ;
        RECT -19.980 -8.360 -19.480 -8.190 ;
        RECT -19.190 -8.360 -18.690 -8.190 ;
        RECT -18.400 -8.360 -17.900 -8.190 ;
        RECT -17.610 -8.360 -17.110 -8.190 ;
        RECT -16.820 -8.360 -16.320 -8.190 ;
        RECT -16.030 -8.360 -15.530 -8.190 ;
        RECT -15.240 -8.360 -14.740 -8.190 ;
        RECT -14.450 -8.360 -13.950 -8.190 ;
        RECT -13.660 -8.360 -13.160 -8.190 ;
        RECT -12.870 -8.360 -12.370 -8.190 ;
        RECT -12.080 -8.360 -11.580 -8.190 ;
        RECT -11.290 -8.360 -10.790 -8.190 ;
        RECT -10.500 -8.360 -10.000 -8.190 ;
        RECT -9.710 -8.360 -9.210 -8.190 ;
        RECT -8.920 -8.360 -8.420 -8.190 ;
        RECT -8.130 -8.360 -7.630 -8.190 ;
        RECT -7.340 -8.360 -6.840 -8.190 ;
        RECT -6.550 -8.360 -6.050 -8.190 ;
        RECT -5.760 -8.360 -5.260 -8.190 ;
        RECT -4.970 -8.360 -4.470 -8.190 ;
        RECT -4.180 -8.360 -3.680 -8.190 ;
        RECT -3.390 -8.360 -2.890 -8.190 ;
        RECT -2.600 -8.360 -2.100 -8.190 ;
        RECT -1.810 -8.360 -1.310 -8.190 ;
        RECT -1.020 -8.360 -0.520 -8.190 ;
        RECT -0.230 -8.360 0.270 -8.190 ;
        RECT 0.560 -8.360 1.060 -8.190 ;
        RECT 1.350 -8.360 1.850 -8.190 ;
        RECT 2.140 -8.360 2.640 -8.190 ;
        RECT 2.930 -8.360 3.430 -8.190 ;
        RECT 3.720 -8.360 4.220 -8.190 ;
        RECT 4.510 -8.360 5.010 -8.190 ;
        RECT 5.300 -8.360 5.800 -8.190 ;
        RECT 6.090 -8.360 6.590 -8.190 ;
        RECT 6.880 -8.360 7.380 -8.190 ;
        RECT 7.670 -8.360 8.170 -8.190 ;
        RECT 8.460 -8.360 8.960 -8.190 ;
        RECT 9.250 -8.360 9.750 -8.190 ;
        RECT 10.040 -8.360 10.540 -8.190 ;
        RECT 10.830 -8.360 11.330 -8.190 ;
        RECT -19.980 -9.910 -19.480 -9.740 ;
        RECT -19.190 -9.910 -18.690 -9.740 ;
        RECT -18.400 -9.910 -17.900 -9.740 ;
        RECT -17.610 -9.910 -17.110 -9.740 ;
        RECT -16.820 -9.910 -16.320 -9.740 ;
        RECT -16.030 -9.910 -15.530 -9.740 ;
        RECT -15.240 -9.910 -14.740 -9.740 ;
        RECT -14.450 -9.910 -13.950 -9.740 ;
        RECT -13.660 -9.910 -13.160 -9.740 ;
        RECT -12.870 -9.910 -12.370 -9.740 ;
        RECT -12.080 -9.910 -11.580 -9.740 ;
        RECT -11.290 -9.910 -10.790 -9.740 ;
        RECT -10.500 -9.910 -10.000 -9.740 ;
        RECT -9.710 -9.910 -9.210 -9.740 ;
        RECT -8.920 -9.910 -8.420 -9.740 ;
        RECT -8.130 -9.910 -7.630 -9.740 ;
        RECT -7.340 -9.910 -6.840 -9.740 ;
        RECT -6.550 -9.910 -6.050 -9.740 ;
        RECT -5.760 -9.910 -5.260 -9.740 ;
        RECT -4.970 -9.910 -4.470 -9.740 ;
        RECT -4.180 -9.910 -3.680 -9.740 ;
        RECT -3.390 -9.910 -2.890 -9.740 ;
        RECT -2.600 -9.910 -2.100 -9.740 ;
        RECT -1.810 -9.910 -1.310 -9.740 ;
        RECT -1.020 -9.910 -0.520 -9.740 ;
        RECT -0.230 -9.910 0.270 -9.740 ;
        RECT 0.560 -9.910 1.060 -9.740 ;
        RECT 1.350 -9.910 1.850 -9.740 ;
        RECT 2.140 -9.910 2.640 -9.740 ;
        RECT 2.930 -9.910 3.430 -9.740 ;
        RECT 3.720 -9.910 4.220 -9.740 ;
        RECT 4.510 -9.910 5.010 -9.740 ;
        RECT 5.300 -9.910 5.800 -9.740 ;
        RECT 6.090 -9.910 6.590 -9.740 ;
        RECT 6.880 -9.910 7.380 -9.740 ;
        RECT 7.670 -9.910 8.170 -9.740 ;
        RECT 8.460 -9.910 8.960 -9.740 ;
        RECT 9.250 -9.910 9.750 -9.740 ;
        RECT 10.040 -9.910 10.540 -9.740 ;
        RECT 10.830 -9.910 11.330 -9.740 ;
        RECT -19.110 -12.180 -16.950 -11.830 ;
        RECT 8.050 -12.180 10.210 -11.830 ;
        RECT -19.110 -13.770 -16.950 -13.420 ;
        RECT 8.050 -13.770 10.210 -13.420 ;
        RECT -19.110 -15.360 -16.950 -15.010 ;
        RECT 8.050 -15.360 10.210 -15.010 ;
        RECT -19.110 -16.950 -16.950 -16.600 ;
      LAYER met1 ;
        RECT -20.855 30.570 12.350 30.890 ;
        RECT -20.855 28.935 -20.535 30.570 ;
        RECT -19.880 30.480 -19.420 30.570 ;
        RECT -19.090 30.480 -18.630 30.570 ;
        RECT -18.300 30.480 -17.840 30.570 ;
        RECT -17.510 30.480 -17.050 30.570 ;
        RECT -16.720 30.480 -16.260 30.570 ;
        RECT -15.930 30.480 -15.470 30.570 ;
        RECT -15.140 30.480 -14.680 30.570 ;
        RECT -14.350 30.480 -13.890 30.570 ;
        RECT -13.560 30.480 -13.100 30.570 ;
        RECT -12.770 30.480 -12.310 30.570 ;
        RECT -11.980 30.480 -11.520 30.570 ;
        RECT -11.190 30.480 -10.730 30.570 ;
        RECT -10.400 30.480 -9.940 30.570 ;
        RECT -9.610 30.480 -9.150 30.570 ;
        RECT -8.820 30.480 -8.360 30.570 ;
        RECT -8.030 30.480 -7.570 30.570 ;
        RECT -7.240 30.480 -6.780 30.570 ;
        RECT -6.450 30.480 -5.990 30.570 ;
        RECT -5.660 30.480 -5.200 30.570 ;
        RECT -4.870 30.480 -4.410 30.570 ;
        RECT -4.080 30.480 -3.620 30.570 ;
        RECT -3.290 30.480 -2.830 30.570 ;
        RECT -2.500 30.480 -2.040 30.570 ;
        RECT -1.710 30.480 -1.250 30.570 ;
        RECT -0.920 30.480 -0.460 30.570 ;
        RECT -0.130 30.480 0.330 30.570 ;
        RECT 0.660 30.480 1.120 30.570 ;
        RECT 1.450 30.480 1.910 30.570 ;
        RECT 2.240 30.480 2.700 30.570 ;
        RECT 3.030 30.480 3.490 30.570 ;
        RECT 3.820 30.480 4.280 30.570 ;
        RECT 4.610 30.480 5.070 30.570 ;
        RECT 5.400 30.480 5.860 30.570 ;
        RECT 6.190 30.480 6.650 30.570 ;
        RECT 6.980 30.480 7.440 30.570 ;
        RECT 7.770 30.480 8.230 30.570 ;
        RECT 8.560 30.480 9.020 30.570 ;
        RECT 9.350 30.480 9.810 30.570 ;
        RECT 10.140 30.480 10.600 30.570 ;
        RECT 10.930 30.480 11.390 30.570 ;
        RECT -19.880 28.935 -19.420 29.070 ;
        RECT -19.090 28.935 -18.630 29.070 ;
        RECT -18.300 28.935 -17.840 29.070 ;
        RECT -17.510 28.935 -17.050 29.070 ;
        RECT -16.720 28.935 -16.260 29.070 ;
        RECT -15.930 28.935 -15.470 29.070 ;
        RECT -15.140 28.935 -14.680 29.070 ;
        RECT -14.350 28.935 -13.890 29.070 ;
        RECT -13.560 28.935 -13.100 29.070 ;
        RECT -12.770 28.935 -12.310 29.070 ;
        RECT -11.980 28.935 -11.520 29.070 ;
        RECT -11.190 28.935 -10.730 29.070 ;
        RECT -10.400 28.935 -9.940 29.070 ;
        RECT -9.610 28.935 -9.150 29.070 ;
        RECT -8.820 28.935 -8.360 29.070 ;
        RECT -8.030 28.935 -7.570 29.070 ;
        RECT -7.240 28.935 -6.780 29.070 ;
        RECT -6.450 28.935 -5.990 29.070 ;
        RECT -5.660 28.935 -5.200 29.070 ;
        RECT -4.870 28.935 -4.410 29.070 ;
        RECT -4.080 28.935 -3.620 29.070 ;
        RECT -3.290 28.935 -2.830 29.070 ;
        RECT -2.500 28.935 -2.040 29.070 ;
        RECT -1.710 28.935 -1.250 29.070 ;
        RECT -0.920 28.935 -0.460 29.070 ;
        RECT -0.130 28.935 0.330 29.070 ;
        RECT 0.660 28.935 1.120 29.070 ;
        RECT 1.450 28.935 1.910 29.070 ;
        RECT 2.240 28.935 2.700 29.070 ;
        RECT 3.030 28.935 3.490 29.070 ;
        RECT 3.820 28.935 4.280 29.070 ;
        RECT 4.610 28.935 5.070 29.070 ;
        RECT 5.400 28.935 5.860 29.070 ;
        RECT 6.190 28.935 6.650 29.070 ;
        RECT 6.980 28.935 7.440 29.070 ;
        RECT 7.770 28.935 8.230 29.070 ;
        RECT 8.560 28.935 9.020 29.070 ;
        RECT 9.350 28.935 9.810 29.070 ;
        RECT 10.140 28.935 10.600 29.070 ;
        RECT 10.930 28.935 11.390 29.070 ;
        RECT 12.030 28.935 12.350 30.570 ;
        RECT -20.855 28.360 12.350 28.935 ;
        RECT -20.855 26.800 -20.535 28.360 ;
        RECT -19.880 28.300 -19.420 28.360 ;
        RECT -19.090 28.300 -18.630 28.360 ;
        RECT -18.300 28.300 -17.840 28.360 ;
        RECT -17.510 28.300 -17.050 28.360 ;
        RECT -16.720 28.300 -16.260 28.360 ;
        RECT -15.930 28.300 -15.470 28.360 ;
        RECT -15.140 28.300 -14.680 28.360 ;
        RECT -14.350 28.300 -13.890 28.360 ;
        RECT -13.560 28.300 -13.100 28.360 ;
        RECT -12.770 28.300 -12.310 28.360 ;
        RECT -11.980 28.300 -11.520 28.360 ;
        RECT -11.190 28.300 -10.730 28.360 ;
        RECT -10.400 28.300 -9.940 28.360 ;
        RECT -9.610 28.300 -9.150 28.360 ;
        RECT -8.820 28.300 -8.360 28.360 ;
        RECT -8.030 28.300 -7.570 28.360 ;
        RECT -7.240 28.300 -6.780 28.360 ;
        RECT -6.450 28.300 -5.990 28.360 ;
        RECT -5.660 28.300 -5.200 28.360 ;
        RECT -4.870 28.300 -4.410 28.360 ;
        RECT -4.080 28.300 -3.620 28.360 ;
        RECT -3.290 28.300 -2.830 28.360 ;
        RECT -2.500 28.300 -2.040 28.360 ;
        RECT -1.710 28.300 -1.250 28.360 ;
        RECT -0.920 28.300 -0.460 28.360 ;
        RECT -0.130 28.300 0.330 28.360 ;
        RECT 0.660 28.300 1.120 28.360 ;
        RECT 1.450 28.300 1.910 28.360 ;
        RECT 2.240 28.300 2.700 28.360 ;
        RECT 3.030 28.300 3.490 28.360 ;
        RECT 3.820 28.300 4.280 28.360 ;
        RECT 4.610 28.300 5.070 28.360 ;
        RECT 5.400 28.300 5.860 28.360 ;
        RECT 6.190 28.300 6.650 28.360 ;
        RECT 6.980 28.300 7.440 28.360 ;
        RECT 7.770 28.300 8.230 28.360 ;
        RECT 8.560 28.300 9.020 28.360 ;
        RECT 9.350 28.300 9.810 28.360 ;
        RECT 10.140 28.300 10.600 28.360 ;
        RECT 10.930 28.300 11.390 28.360 ;
        RECT -19.880 26.800 -19.420 26.890 ;
        RECT -19.090 26.800 -18.630 26.890 ;
        RECT -18.300 26.800 -17.840 26.890 ;
        RECT -17.510 26.800 -17.050 26.890 ;
        RECT -16.720 26.800 -16.260 26.890 ;
        RECT -15.930 26.800 -15.470 26.890 ;
        RECT -15.140 26.800 -14.680 26.890 ;
        RECT -14.350 26.800 -13.890 26.890 ;
        RECT -13.560 26.800 -13.100 26.890 ;
        RECT -12.770 26.800 -12.310 26.890 ;
        RECT -11.980 26.800 -11.520 26.890 ;
        RECT -11.190 26.800 -10.730 26.890 ;
        RECT -10.400 26.800 -9.940 26.890 ;
        RECT -9.610 26.800 -9.150 26.890 ;
        RECT -8.820 26.800 -8.360 26.890 ;
        RECT -8.030 26.800 -7.570 26.890 ;
        RECT -7.240 26.800 -6.780 26.890 ;
        RECT -6.450 26.800 -5.990 26.890 ;
        RECT -5.660 26.800 -5.200 26.890 ;
        RECT -4.870 26.800 -4.410 26.890 ;
        RECT -4.080 26.800 -3.620 26.890 ;
        RECT -3.290 26.800 -2.830 26.890 ;
        RECT -2.500 26.800 -2.040 26.890 ;
        RECT -1.710 26.800 -1.250 26.890 ;
        RECT -0.920 26.800 -0.460 26.890 ;
        RECT -0.130 26.800 0.330 26.890 ;
        RECT 0.660 26.800 1.120 26.890 ;
        RECT 1.450 26.800 1.910 26.890 ;
        RECT 2.240 26.800 2.700 26.890 ;
        RECT 3.030 26.800 3.490 26.890 ;
        RECT 3.820 26.800 4.280 26.890 ;
        RECT 4.610 26.800 5.070 26.890 ;
        RECT 5.400 26.800 5.860 26.890 ;
        RECT 6.190 26.800 6.650 26.890 ;
        RECT 6.980 26.800 7.440 26.890 ;
        RECT 7.770 26.800 8.230 26.890 ;
        RECT 8.560 26.800 9.020 26.890 ;
        RECT 9.350 26.800 9.810 26.890 ;
        RECT 10.140 26.800 10.600 26.890 ;
        RECT 10.930 26.800 11.390 26.890 ;
        RECT 12.030 26.800 12.350 28.360 ;
        RECT -20.855 26.225 12.350 26.800 ;
        RECT -20.855 24.585 -20.535 26.225 ;
        RECT -19.880 26.120 -19.420 26.225 ;
        RECT -19.090 26.120 -18.630 26.225 ;
        RECT -18.300 26.120 -17.840 26.225 ;
        RECT -17.510 26.120 -17.050 26.225 ;
        RECT -16.720 26.120 -16.260 26.225 ;
        RECT -15.930 26.120 -15.470 26.225 ;
        RECT -15.140 26.120 -14.680 26.225 ;
        RECT -14.350 26.120 -13.890 26.225 ;
        RECT -13.560 26.120 -13.100 26.225 ;
        RECT -12.770 26.120 -12.310 26.225 ;
        RECT -11.980 26.120 -11.520 26.225 ;
        RECT -11.190 26.120 -10.730 26.225 ;
        RECT -10.400 26.120 -9.940 26.225 ;
        RECT -9.610 26.120 -9.150 26.225 ;
        RECT -8.820 26.120 -8.360 26.225 ;
        RECT -8.030 26.120 -7.570 26.225 ;
        RECT -7.240 26.120 -6.780 26.225 ;
        RECT -6.450 26.120 -5.990 26.225 ;
        RECT -5.660 26.120 -5.200 26.225 ;
        RECT -4.870 26.120 -4.410 26.225 ;
        RECT -4.080 26.120 -3.620 26.225 ;
        RECT -3.290 26.120 -2.830 26.225 ;
        RECT -2.500 26.120 -2.040 26.225 ;
        RECT -1.710 26.120 -1.250 26.225 ;
        RECT -0.920 26.120 -0.460 26.225 ;
        RECT -0.130 26.120 0.330 26.225 ;
        RECT 0.660 26.120 1.120 26.225 ;
        RECT 1.450 26.120 1.910 26.225 ;
        RECT 2.240 26.120 2.700 26.225 ;
        RECT 3.030 26.120 3.490 26.225 ;
        RECT 3.820 26.120 4.280 26.225 ;
        RECT 4.610 26.120 5.070 26.225 ;
        RECT 5.400 26.120 5.860 26.225 ;
        RECT 6.190 26.120 6.650 26.225 ;
        RECT 6.980 26.120 7.440 26.225 ;
        RECT 7.770 26.120 8.230 26.225 ;
        RECT 8.560 26.120 9.020 26.225 ;
        RECT 9.350 26.120 9.810 26.225 ;
        RECT 10.140 26.120 10.600 26.225 ;
        RECT 10.930 26.120 11.390 26.225 ;
        RECT -19.880 24.585 -19.420 24.710 ;
        RECT -19.090 24.585 -18.630 24.710 ;
        RECT -18.300 24.585 -17.840 24.710 ;
        RECT -17.510 24.585 -17.050 24.710 ;
        RECT -16.720 24.585 -16.260 24.710 ;
        RECT -15.930 24.585 -15.470 24.710 ;
        RECT -15.140 24.585 -14.680 24.710 ;
        RECT -14.350 24.585 -13.890 24.710 ;
        RECT -13.560 24.585 -13.100 24.710 ;
        RECT -12.770 24.585 -12.310 24.710 ;
        RECT -11.980 24.585 -11.520 24.710 ;
        RECT -11.190 24.585 -10.730 24.710 ;
        RECT -10.400 24.585 -9.940 24.710 ;
        RECT -9.610 24.585 -9.150 24.710 ;
        RECT -8.820 24.585 -8.360 24.710 ;
        RECT -8.030 24.585 -7.570 24.710 ;
        RECT -7.240 24.585 -6.780 24.710 ;
        RECT -6.450 24.585 -5.990 24.710 ;
        RECT -5.660 24.585 -5.200 24.710 ;
        RECT -4.870 24.585 -4.410 24.710 ;
        RECT -4.080 24.585 -3.620 24.710 ;
        RECT -3.290 24.585 -2.830 24.710 ;
        RECT -2.500 24.585 -2.040 24.710 ;
        RECT -1.710 24.585 -1.250 24.710 ;
        RECT -0.920 24.585 -0.460 24.710 ;
        RECT -0.130 24.585 0.330 24.710 ;
        RECT 0.660 24.585 1.120 24.710 ;
        RECT 1.450 24.585 1.910 24.710 ;
        RECT 2.240 24.585 2.700 24.710 ;
        RECT 3.030 24.585 3.490 24.710 ;
        RECT 3.820 24.585 4.280 24.710 ;
        RECT 4.610 24.585 5.070 24.710 ;
        RECT 5.400 24.585 5.860 24.710 ;
        RECT 6.190 24.585 6.650 24.710 ;
        RECT 6.980 24.585 7.440 24.710 ;
        RECT 7.770 24.585 8.230 24.710 ;
        RECT 8.560 24.585 9.020 24.710 ;
        RECT 9.350 24.585 9.810 24.710 ;
        RECT 10.140 24.585 10.600 24.710 ;
        RECT 10.930 24.585 11.390 24.710 ;
        RECT 12.030 24.585 12.350 26.225 ;
        RECT -20.855 24.010 12.350 24.585 ;
        RECT -20.855 22.420 -20.535 24.010 ;
        RECT -19.880 23.940 -19.420 24.010 ;
        RECT -19.090 23.940 -18.630 24.010 ;
        RECT -18.300 23.940 -17.840 24.010 ;
        RECT -17.510 23.940 -17.050 24.010 ;
        RECT -16.720 23.940 -16.260 24.010 ;
        RECT -15.930 23.940 -15.470 24.010 ;
        RECT -15.140 23.940 -14.680 24.010 ;
        RECT -14.350 23.940 -13.890 24.010 ;
        RECT -13.560 23.940 -13.100 24.010 ;
        RECT -12.770 23.940 -12.310 24.010 ;
        RECT -11.980 23.940 -11.520 24.010 ;
        RECT -11.190 23.940 -10.730 24.010 ;
        RECT -10.400 23.940 -9.940 24.010 ;
        RECT -9.610 23.940 -9.150 24.010 ;
        RECT -8.820 23.940 -8.360 24.010 ;
        RECT -8.030 23.940 -7.570 24.010 ;
        RECT -7.240 23.940 -6.780 24.010 ;
        RECT -6.450 23.940 -5.990 24.010 ;
        RECT -5.660 23.940 -5.200 24.010 ;
        RECT -4.870 23.940 -4.410 24.010 ;
        RECT -4.080 23.940 -3.620 24.010 ;
        RECT -3.290 23.940 -2.830 24.010 ;
        RECT -2.500 23.940 -2.040 24.010 ;
        RECT -1.710 23.940 -1.250 24.010 ;
        RECT -0.920 23.940 -0.460 24.010 ;
        RECT -0.130 23.940 0.330 24.010 ;
        RECT 0.660 23.940 1.120 24.010 ;
        RECT 1.450 23.940 1.910 24.010 ;
        RECT 2.240 23.940 2.700 24.010 ;
        RECT 3.030 23.940 3.490 24.010 ;
        RECT 3.820 23.940 4.280 24.010 ;
        RECT 4.610 23.940 5.070 24.010 ;
        RECT 5.400 23.940 5.860 24.010 ;
        RECT 6.190 23.940 6.650 24.010 ;
        RECT 6.980 23.940 7.440 24.010 ;
        RECT 7.770 23.940 8.230 24.010 ;
        RECT 8.560 23.940 9.020 24.010 ;
        RECT 9.350 23.940 9.810 24.010 ;
        RECT 10.140 23.940 10.600 24.010 ;
        RECT 10.930 23.940 11.390 24.010 ;
        RECT -19.880 22.420 -19.420 22.530 ;
        RECT -19.090 22.420 -18.630 22.530 ;
        RECT -18.300 22.420 -17.840 22.530 ;
        RECT -17.510 22.420 -17.050 22.530 ;
        RECT -16.720 22.420 -16.260 22.530 ;
        RECT -15.930 22.420 -15.470 22.530 ;
        RECT -15.140 22.420 -14.680 22.530 ;
        RECT -14.350 22.420 -13.890 22.530 ;
        RECT -13.560 22.420 -13.100 22.530 ;
        RECT -12.770 22.420 -12.310 22.530 ;
        RECT -11.980 22.420 -11.520 22.530 ;
        RECT -11.190 22.420 -10.730 22.530 ;
        RECT -10.400 22.420 -9.940 22.530 ;
        RECT -9.610 22.420 -9.150 22.530 ;
        RECT -8.820 22.420 -8.360 22.530 ;
        RECT -8.030 22.420 -7.570 22.530 ;
        RECT -7.240 22.420 -6.780 22.530 ;
        RECT -6.450 22.420 -5.990 22.530 ;
        RECT -5.660 22.420 -5.200 22.530 ;
        RECT -4.870 22.420 -4.410 22.530 ;
        RECT -4.080 22.420 -3.620 22.530 ;
        RECT -3.290 22.420 -2.830 22.530 ;
        RECT -2.500 22.420 -2.040 22.530 ;
        RECT -1.710 22.420 -1.250 22.530 ;
        RECT -0.920 22.420 -0.460 22.530 ;
        RECT -0.130 22.420 0.330 22.530 ;
        RECT 0.660 22.420 1.120 22.530 ;
        RECT 1.450 22.420 1.910 22.530 ;
        RECT 2.240 22.420 2.700 22.530 ;
        RECT 3.030 22.420 3.490 22.530 ;
        RECT 3.820 22.420 4.280 22.530 ;
        RECT 4.610 22.420 5.070 22.530 ;
        RECT 5.400 22.420 5.860 22.530 ;
        RECT 6.190 22.420 6.650 22.530 ;
        RECT 6.980 22.420 7.440 22.530 ;
        RECT 7.770 22.420 8.230 22.530 ;
        RECT 8.560 22.420 9.020 22.530 ;
        RECT 9.350 22.420 9.810 22.530 ;
        RECT 10.140 22.420 10.600 22.530 ;
        RECT 10.930 22.420 11.390 22.530 ;
        RECT 12.030 22.420 12.350 24.010 ;
        RECT -20.855 21.845 12.350 22.420 ;
        RECT -20.855 20.355 -20.535 21.845 ;
        RECT -19.880 21.760 -19.420 21.845 ;
        RECT -19.090 21.760 -18.630 21.845 ;
        RECT -18.300 21.760 -17.840 21.845 ;
        RECT -17.510 21.760 -17.050 21.845 ;
        RECT -16.720 21.760 -16.260 21.845 ;
        RECT -15.930 21.760 -15.470 21.845 ;
        RECT -15.140 21.760 -14.680 21.845 ;
        RECT -14.350 21.760 -13.890 21.845 ;
        RECT -13.560 21.760 -13.100 21.845 ;
        RECT -12.770 21.760 -12.310 21.845 ;
        RECT -11.980 21.760 -11.520 21.845 ;
        RECT -11.190 21.760 -10.730 21.845 ;
        RECT -10.400 21.760 -9.940 21.845 ;
        RECT -9.610 21.760 -9.150 21.845 ;
        RECT -8.820 21.760 -8.360 21.845 ;
        RECT -8.030 21.760 -7.570 21.845 ;
        RECT -7.240 21.760 -6.780 21.845 ;
        RECT -6.450 21.760 -5.990 21.845 ;
        RECT -5.660 21.760 -5.200 21.845 ;
        RECT -4.870 21.760 -4.410 21.845 ;
        RECT -4.080 21.760 -3.620 21.845 ;
        RECT -3.290 21.760 -2.830 21.845 ;
        RECT -2.500 21.760 -2.040 21.845 ;
        RECT -1.710 21.760 -1.250 21.845 ;
        RECT -0.920 21.760 -0.460 21.845 ;
        RECT -0.130 21.760 0.330 21.845 ;
        RECT 0.660 21.760 1.120 21.845 ;
        RECT 1.450 21.760 1.910 21.845 ;
        RECT 2.240 21.760 2.700 21.845 ;
        RECT 3.030 21.760 3.490 21.845 ;
        RECT 3.820 21.760 4.280 21.845 ;
        RECT 4.610 21.760 5.070 21.845 ;
        RECT 5.400 21.760 5.860 21.845 ;
        RECT 6.190 21.760 6.650 21.845 ;
        RECT 6.980 21.760 7.440 21.845 ;
        RECT 7.770 21.760 8.230 21.845 ;
        RECT 8.560 21.760 9.020 21.845 ;
        RECT 9.350 21.760 9.810 21.845 ;
        RECT 10.140 21.760 10.600 21.845 ;
        RECT 10.930 21.760 11.390 21.845 ;
        RECT -21.455 20.330 -20.535 20.355 ;
        RECT -19.880 20.330 -19.420 20.350 ;
        RECT -19.090 20.330 -18.630 20.350 ;
        RECT -18.300 20.330 -17.840 20.350 ;
        RECT -17.510 20.330 -17.050 20.350 ;
        RECT -16.720 20.330 -16.260 20.350 ;
        RECT -15.930 20.330 -15.470 20.350 ;
        RECT -15.140 20.330 -14.680 20.350 ;
        RECT -14.350 20.330 -13.890 20.350 ;
        RECT -13.560 20.330 -13.100 20.350 ;
        RECT -12.770 20.330 -12.310 20.350 ;
        RECT -11.980 20.330 -11.520 20.350 ;
        RECT -11.190 20.330 -10.730 20.350 ;
        RECT -10.400 20.330 -9.940 20.350 ;
        RECT -9.610 20.330 -9.150 20.350 ;
        RECT -8.820 20.330 -8.360 20.350 ;
        RECT -8.030 20.330 -7.570 20.350 ;
        RECT -7.240 20.330 -6.780 20.350 ;
        RECT -6.450 20.330 -5.990 20.350 ;
        RECT -5.660 20.330 -5.200 20.350 ;
        RECT -4.870 20.330 -4.410 20.350 ;
        RECT -4.080 20.330 -3.620 20.350 ;
        RECT -3.290 20.330 -2.830 20.350 ;
        RECT -2.500 20.330 -2.040 20.350 ;
        RECT -1.710 20.330 -1.250 20.350 ;
        RECT -0.920 20.330 -0.460 20.350 ;
        RECT -0.130 20.330 0.330 20.350 ;
        RECT 0.660 20.330 1.120 20.350 ;
        RECT 1.450 20.330 1.910 20.350 ;
        RECT 2.240 20.330 2.700 20.350 ;
        RECT 3.030 20.330 3.490 20.350 ;
        RECT 3.820 20.330 4.280 20.350 ;
        RECT 4.610 20.330 5.070 20.350 ;
        RECT 5.400 20.330 5.860 20.350 ;
        RECT 6.190 20.330 6.650 20.350 ;
        RECT 6.980 20.330 7.440 20.350 ;
        RECT 7.770 20.330 8.230 20.350 ;
        RECT 8.560 20.330 9.020 20.350 ;
        RECT 9.350 20.330 9.810 20.350 ;
        RECT 10.140 20.330 10.600 20.350 ;
        RECT 10.930 20.330 11.390 20.350 ;
        RECT 12.030 20.330 12.350 21.845 ;
        RECT -21.455 20.010 12.350 20.330 ;
        RECT -21.455 7.915 -21.135 20.010 ;
        RECT -20.870 18.785 12.380 19.105 ;
        RECT -20.870 17.200 -20.550 18.785 ;
        RECT -19.880 18.740 -19.420 18.785 ;
        RECT -19.090 18.740 -18.630 18.785 ;
        RECT -18.300 18.740 -17.840 18.785 ;
        RECT -17.510 18.740 -17.050 18.785 ;
        RECT -16.720 18.740 -16.260 18.785 ;
        RECT -15.930 18.740 -15.470 18.785 ;
        RECT -15.140 18.740 -14.680 18.785 ;
        RECT -14.350 18.740 -13.890 18.785 ;
        RECT -13.560 18.740 -13.100 18.785 ;
        RECT -12.770 18.740 -12.310 18.785 ;
        RECT -11.980 18.740 -11.520 18.785 ;
        RECT -11.190 18.740 -10.730 18.785 ;
        RECT -10.400 18.740 -9.940 18.785 ;
        RECT -9.610 18.740 -9.150 18.785 ;
        RECT -8.820 18.740 -8.360 18.785 ;
        RECT -8.030 18.740 -7.570 18.785 ;
        RECT -7.240 18.740 -6.780 18.785 ;
        RECT -6.450 18.740 -5.990 18.785 ;
        RECT -5.660 18.740 -5.200 18.785 ;
        RECT -4.870 18.740 -4.410 18.785 ;
        RECT -4.080 18.740 -3.620 18.785 ;
        RECT -3.290 18.740 -2.830 18.785 ;
        RECT -2.500 18.740 -2.040 18.785 ;
        RECT -1.710 18.740 -1.250 18.785 ;
        RECT -0.920 18.740 -0.460 18.785 ;
        RECT -0.130 18.740 0.330 18.785 ;
        RECT 0.660 18.740 1.120 18.785 ;
        RECT 1.450 18.740 1.910 18.785 ;
        RECT 2.240 18.740 2.700 18.785 ;
        RECT 3.030 18.740 3.490 18.785 ;
        RECT 3.820 18.740 4.280 18.785 ;
        RECT 4.610 18.740 5.070 18.785 ;
        RECT 5.400 18.740 5.860 18.785 ;
        RECT 6.190 18.740 6.650 18.785 ;
        RECT 6.980 18.740 7.440 18.785 ;
        RECT 7.770 18.740 8.230 18.785 ;
        RECT 8.560 18.740 9.020 18.785 ;
        RECT 9.350 18.740 9.810 18.785 ;
        RECT 10.140 18.740 10.600 18.785 ;
        RECT 10.930 18.740 11.390 18.785 ;
        RECT -19.880 17.200 -19.420 17.330 ;
        RECT -19.090 17.200 -18.630 17.330 ;
        RECT -18.300 17.200 -17.840 17.330 ;
        RECT -17.510 17.200 -17.050 17.330 ;
        RECT -16.720 17.200 -16.260 17.330 ;
        RECT -15.930 17.200 -15.470 17.330 ;
        RECT -15.140 17.200 -14.680 17.330 ;
        RECT -14.350 17.200 -13.890 17.330 ;
        RECT -13.560 17.200 -13.100 17.330 ;
        RECT -12.770 17.200 -12.310 17.330 ;
        RECT -11.980 17.200 -11.520 17.330 ;
        RECT -11.190 17.200 -10.730 17.330 ;
        RECT -10.400 17.200 -9.940 17.330 ;
        RECT -9.610 17.200 -9.150 17.330 ;
        RECT -8.820 17.200 -8.360 17.330 ;
        RECT -8.030 17.200 -7.570 17.330 ;
        RECT -7.240 17.200 -6.780 17.330 ;
        RECT -6.450 17.200 -5.990 17.330 ;
        RECT -5.660 17.200 -5.200 17.330 ;
        RECT -4.870 17.200 -4.410 17.330 ;
        RECT -4.080 17.200 -3.620 17.330 ;
        RECT -3.290 17.200 -2.830 17.330 ;
        RECT -2.500 17.200 -2.040 17.330 ;
        RECT -1.710 17.200 -1.250 17.330 ;
        RECT -0.920 17.200 -0.460 17.330 ;
        RECT -0.130 17.200 0.330 17.330 ;
        RECT 0.660 17.200 1.120 17.330 ;
        RECT 1.450 17.200 1.910 17.330 ;
        RECT 2.240 17.200 2.700 17.330 ;
        RECT 3.030 17.200 3.490 17.330 ;
        RECT 3.820 17.200 4.280 17.330 ;
        RECT 4.610 17.200 5.070 17.330 ;
        RECT 5.400 17.200 5.860 17.330 ;
        RECT 6.190 17.200 6.650 17.330 ;
        RECT 6.980 17.200 7.440 17.330 ;
        RECT 7.770 17.200 8.230 17.330 ;
        RECT 8.560 17.200 9.020 17.330 ;
        RECT 9.350 17.200 9.810 17.330 ;
        RECT 10.140 17.200 10.600 17.330 ;
        RECT 10.930 17.200 11.390 17.330 ;
        RECT 12.060 17.200 12.380 18.785 ;
        RECT -20.870 16.625 12.380 17.200 ;
        RECT -20.870 15.010 -20.550 16.625 ;
        RECT -19.880 16.560 -19.420 16.625 ;
        RECT -19.090 16.560 -18.630 16.625 ;
        RECT -18.300 16.560 -17.840 16.625 ;
        RECT -17.510 16.560 -17.050 16.625 ;
        RECT -16.720 16.560 -16.260 16.625 ;
        RECT -15.930 16.560 -15.470 16.625 ;
        RECT -15.140 16.560 -14.680 16.625 ;
        RECT -14.350 16.560 -13.890 16.625 ;
        RECT -13.560 16.560 -13.100 16.625 ;
        RECT -12.770 16.560 -12.310 16.625 ;
        RECT -11.980 16.560 -11.520 16.625 ;
        RECT -11.190 16.560 -10.730 16.625 ;
        RECT -10.400 16.560 -9.940 16.625 ;
        RECT -9.610 16.560 -9.150 16.625 ;
        RECT -8.820 16.560 -8.360 16.625 ;
        RECT -8.030 16.560 -7.570 16.625 ;
        RECT -7.240 16.560 -6.780 16.625 ;
        RECT -6.450 16.560 -5.990 16.625 ;
        RECT -5.660 16.560 -5.200 16.625 ;
        RECT -4.870 16.560 -4.410 16.625 ;
        RECT -4.080 16.560 -3.620 16.625 ;
        RECT -3.290 16.560 -2.830 16.625 ;
        RECT -2.500 16.560 -2.040 16.625 ;
        RECT -1.710 16.560 -1.250 16.625 ;
        RECT -0.920 16.560 -0.460 16.625 ;
        RECT -0.130 16.560 0.330 16.625 ;
        RECT 0.660 16.560 1.120 16.625 ;
        RECT 1.450 16.560 1.910 16.625 ;
        RECT 2.240 16.560 2.700 16.625 ;
        RECT 3.030 16.560 3.490 16.625 ;
        RECT 3.820 16.560 4.280 16.625 ;
        RECT 4.610 16.560 5.070 16.625 ;
        RECT 5.400 16.560 5.860 16.625 ;
        RECT 6.190 16.560 6.650 16.625 ;
        RECT 6.980 16.560 7.440 16.625 ;
        RECT 7.770 16.560 8.230 16.625 ;
        RECT 8.560 16.560 9.020 16.625 ;
        RECT 9.350 16.560 9.810 16.625 ;
        RECT 10.140 16.560 10.600 16.625 ;
        RECT 10.930 16.560 11.390 16.625 ;
        RECT -19.880 15.010 -19.420 15.150 ;
        RECT -19.090 15.010 -18.630 15.150 ;
        RECT -18.300 15.010 -17.840 15.150 ;
        RECT -17.510 15.010 -17.050 15.150 ;
        RECT -16.720 15.010 -16.260 15.150 ;
        RECT -15.930 15.010 -15.470 15.150 ;
        RECT -15.140 15.010 -14.680 15.150 ;
        RECT -14.350 15.010 -13.890 15.150 ;
        RECT -13.560 15.010 -13.100 15.150 ;
        RECT -12.770 15.010 -12.310 15.150 ;
        RECT -11.980 15.010 -11.520 15.150 ;
        RECT -11.190 15.010 -10.730 15.150 ;
        RECT -10.400 15.010 -9.940 15.150 ;
        RECT -9.610 15.010 -9.150 15.150 ;
        RECT -8.820 15.010 -8.360 15.150 ;
        RECT -8.030 15.010 -7.570 15.150 ;
        RECT -7.240 15.010 -6.780 15.150 ;
        RECT -6.450 15.010 -5.990 15.150 ;
        RECT -5.660 15.010 -5.200 15.150 ;
        RECT -4.870 15.010 -4.410 15.150 ;
        RECT -4.080 15.010 -3.620 15.150 ;
        RECT -3.290 15.010 -2.830 15.150 ;
        RECT -2.500 15.010 -2.040 15.150 ;
        RECT -1.710 15.010 -1.250 15.150 ;
        RECT -0.920 15.010 -0.460 15.150 ;
        RECT -0.130 15.010 0.330 15.150 ;
        RECT 0.660 15.010 1.120 15.150 ;
        RECT 1.450 15.010 1.910 15.150 ;
        RECT 2.240 15.010 2.700 15.150 ;
        RECT 3.030 15.010 3.490 15.150 ;
        RECT 3.820 15.010 4.280 15.150 ;
        RECT 4.610 15.010 5.070 15.150 ;
        RECT 5.400 15.010 5.860 15.150 ;
        RECT 6.190 15.010 6.650 15.150 ;
        RECT 6.980 15.010 7.440 15.150 ;
        RECT 7.770 15.010 8.230 15.150 ;
        RECT 8.560 15.010 9.020 15.150 ;
        RECT 9.350 15.010 9.810 15.150 ;
        RECT 10.140 15.010 10.600 15.150 ;
        RECT 10.930 15.010 11.390 15.150 ;
        RECT 12.060 15.010 12.380 16.625 ;
        RECT -20.870 14.435 12.380 15.010 ;
        RECT -20.870 12.850 -20.550 14.435 ;
        RECT -19.880 14.380 -19.420 14.435 ;
        RECT -19.090 14.380 -18.630 14.435 ;
        RECT -18.300 14.380 -17.840 14.435 ;
        RECT -17.510 14.380 -17.050 14.435 ;
        RECT -16.720 14.380 -16.260 14.435 ;
        RECT -15.930 14.380 -15.470 14.435 ;
        RECT -15.140 14.380 -14.680 14.435 ;
        RECT -14.350 14.380 -13.890 14.435 ;
        RECT -13.560 14.380 -13.100 14.435 ;
        RECT -12.770 14.380 -12.310 14.435 ;
        RECT -11.980 14.380 -11.520 14.435 ;
        RECT -11.190 14.380 -10.730 14.435 ;
        RECT -10.400 14.380 -9.940 14.435 ;
        RECT -9.610 14.380 -9.150 14.435 ;
        RECT -8.820 14.380 -8.360 14.435 ;
        RECT -8.030 14.380 -7.570 14.435 ;
        RECT -7.240 14.380 -6.780 14.435 ;
        RECT -6.450 14.380 -5.990 14.435 ;
        RECT -5.660 14.380 -5.200 14.435 ;
        RECT -4.870 14.380 -4.410 14.435 ;
        RECT -4.080 14.380 -3.620 14.435 ;
        RECT -3.290 14.380 -2.830 14.435 ;
        RECT -2.500 14.380 -2.040 14.435 ;
        RECT -1.710 14.380 -1.250 14.435 ;
        RECT -0.920 14.380 -0.460 14.435 ;
        RECT -0.130 14.380 0.330 14.435 ;
        RECT 0.660 14.380 1.120 14.435 ;
        RECT 1.450 14.380 1.910 14.435 ;
        RECT 2.240 14.380 2.700 14.435 ;
        RECT 3.030 14.380 3.490 14.435 ;
        RECT 3.820 14.380 4.280 14.435 ;
        RECT 4.610 14.380 5.070 14.435 ;
        RECT 5.400 14.380 5.860 14.435 ;
        RECT 6.190 14.380 6.650 14.435 ;
        RECT 6.980 14.380 7.440 14.435 ;
        RECT 7.770 14.380 8.230 14.435 ;
        RECT 8.560 14.380 9.020 14.435 ;
        RECT 9.350 14.380 9.810 14.435 ;
        RECT 10.140 14.380 10.600 14.435 ;
        RECT 10.930 14.380 11.390 14.435 ;
        RECT -19.880 12.850 -19.420 12.970 ;
        RECT -19.090 12.850 -18.630 12.970 ;
        RECT -18.300 12.850 -17.840 12.970 ;
        RECT -17.510 12.850 -17.050 12.970 ;
        RECT -16.720 12.850 -16.260 12.970 ;
        RECT -15.930 12.850 -15.470 12.970 ;
        RECT -15.140 12.850 -14.680 12.970 ;
        RECT -14.350 12.850 -13.890 12.970 ;
        RECT -13.560 12.850 -13.100 12.970 ;
        RECT -12.770 12.850 -12.310 12.970 ;
        RECT -11.980 12.850 -11.520 12.970 ;
        RECT -11.190 12.850 -10.730 12.970 ;
        RECT -10.400 12.850 -9.940 12.970 ;
        RECT -9.610 12.850 -9.150 12.970 ;
        RECT -8.820 12.850 -8.360 12.970 ;
        RECT -8.030 12.850 -7.570 12.970 ;
        RECT -7.240 12.850 -6.780 12.970 ;
        RECT -6.450 12.850 -5.990 12.970 ;
        RECT -5.660 12.850 -5.200 12.970 ;
        RECT -4.870 12.850 -4.410 12.970 ;
        RECT -4.080 12.850 -3.620 12.970 ;
        RECT -3.290 12.850 -2.830 12.970 ;
        RECT -2.500 12.850 -2.040 12.970 ;
        RECT -1.710 12.850 -1.250 12.970 ;
        RECT -0.920 12.850 -0.460 12.970 ;
        RECT -0.130 12.850 0.330 12.970 ;
        RECT 0.660 12.850 1.120 12.970 ;
        RECT 1.450 12.850 1.910 12.970 ;
        RECT 2.240 12.850 2.700 12.970 ;
        RECT 3.030 12.850 3.490 12.970 ;
        RECT 3.820 12.850 4.280 12.970 ;
        RECT 4.610 12.850 5.070 12.970 ;
        RECT 5.400 12.850 5.860 12.970 ;
        RECT 6.190 12.850 6.650 12.970 ;
        RECT 6.980 12.850 7.440 12.970 ;
        RECT 7.770 12.850 8.230 12.970 ;
        RECT 8.560 12.850 9.020 12.970 ;
        RECT 9.350 12.850 9.810 12.970 ;
        RECT 10.140 12.850 10.600 12.970 ;
        RECT 10.930 12.850 11.390 12.970 ;
        RECT 12.060 12.850 12.380 14.435 ;
        RECT -20.870 12.275 12.380 12.850 ;
        RECT -20.870 10.675 -20.550 12.275 ;
        RECT -19.880 12.200 -19.420 12.275 ;
        RECT -19.090 12.200 -18.630 12.275 ;
        RECT -18.300 12.200 -17.840 12.275 ;
        RECT -17.510 12.200 -17.050 12.275 ;
        RECT -16.720 12.200 -16.260 12.275 ;
        RECT -15.930 12.200 -15.470 12.275 ;
        RECT -15.140 12.200 -14.680 12.275 ;
        RECT -14.350 12.200 -13.890 12.275 ;
        RECT -13.560 12.200 -13.100 12.275 ;
        RECT -12.770 12.200 -12.310 12.275 ;
        RECT -11.980 12.200 -11.520 12.275 ;
        RECT -11.190 12.200 -10.730 12.275 ;
        RECT -10.400 12.200 -9.940 12.275 ;
        RECT -9.610 12.200 -9.150 12.275 ;
        RECT -8.820 12.200 -8.360 12.275 ;
        RECT -8.030 12.200 -7.570 12.275 ;
        RECT -7.240 12.200 -6.780 12.275 ;
        RECT -6.450 12.200 -5.990 12.275 ;
        RECT -5.660 12.200 -5.200 12.275 ;
        RECT -4.870 12.200 -4.410 12.275 ;
        RECT -4.080 12.200 -3.620 12.275 ;
        RECT -3.290 12.200 -2.830 12.275 ;
        RECT -2.500 12.200 -2.040 12.275 ;
        RECT -1.710 12.200 -1.250 12.275 ;
        RECT -0.920 12.200 -0.460 12.275 ;
        RECT -0.130 12.200 0.330 12.275 ;
        RECT 0.660 12.200 1.120 12.275 ;
        RECT 1.450 12.200 1.910 12.275 ;
        RECT 2.240 12.200 2.700 12.275 ;
        RECT 3.030 12.200 3.490 12.275 ;
        RECT 3.820 12.200 4.280 12.275 ;
        RECT 4.610 12.200 5.070 12.275 ;
        RECT 5.400 12.200 5.860 12.275 ;
        RECT 6.190 12.200 6.650 12.275 ;
        RECT 6.980 12.200 7.440 12.275 ;
        RECT 7.770 12.200 8.230 12.275 ;
        RECT 8.560 12.200 9.020 12.275 ;
        RECT 9.350 12.200 9.810 12.275 ;
        RECT 10.140 12.200 10.600 12.275 ;
        RECT 10.930 12.200 11.390 12.275 ;
        RECT -19.880 10.675 -19.420 10.790 ;
        RECT -19.090 10.675 -18.630 10.790 ;
        RECT -18.300 10.675 -17.840 10.790 ;
        RECT -17.510 10.675 -17.050 10.790 ;
        RECT -16.720 10.675 -16.260 10.790 ;
        RECT -15.930 10.675 -15.470 10.790 ;
        RECT -15.140 10.675 -14.680 10.790 ;
        RECT -14.350 10.675 -13.890 10.790 ;
        RECT -13.560 10.675 -13.100 10.790 ;
        RECT -12.770 10.675 -12.310 10.790 ;
        RECT -11.980 10.675 -11.520 10.790 ;
        RECT -11.190 10.675 -10.730 10.790 ;
        RECT -10.400 10.675 -9.940 10.790 ;
        RECT -9.610 10.675 -9.150 10.790 ;
        RECT -8.820 10.675 -8.360 10.790 ;
        RECT -8.030 10.675 -7.570 10.790 ;
        RECT -7.240 10.675 -6.780 10.790 ;
        RECT -6.450 10.675 -5.990 10.790 ;
        RECT -5.660 10.675 -5.200 10.790 ;
        RECT -4.870 10.675 -4.410 10.790 ;
        RECT -4.080 10.675 -3.620 10.790 ;
        RECT -3.290 10.675 -2.830 10.790 ;
        RECT -2.500 10.675 -2.040 10.790 ;
        RECT -1.710 10.675 -1.250 10.790 ;
        RECT -0.920 10.675 -0.460 10.790 ;
        RECT -0.130 10.675 0.330 10.790 ;
        RECT 0.660 10.675 1.120 10.790 ;
        RECT 1.450 10.675 1.910 10.790 ;
        RECT 2.240 10.675 2.700 10.790 ;
        RECT 3.030 10.675 3.490 10.790 ;
        RECT 3.820 10.675 4.280 10.790 ;
        RECT 4.610 10.675 5.070 10.790 ;
        RECT 5.400 10.675 5.860 10.790 ;
        RECT 6.190 10.675 6.650 10.790 ;
        RECT 6.980 10.675 7.440 10.790 ;
        RECT 7.770 10.675 8.230 10.790 ;
        RECT 8.560 10.675 9.020 10.790 ;
        RECT 9.350 10.675 9.810 10.790 ;
        RECT 10.140 10.675 10.600 10.790 ;
        RECT 10.930 10.675 11.390 10.790 ;
        RECT 12.060 10.675 12.380 12.275 ;
        RECT -20.870 10.200 12.380 10.675 ;
        RECT -20.870 8.565 -20.550 10.200 ;
        RECT -19.880 10.020 -19.420 10.200 ;
        RECT -19.090 10.020 -18.630 10.200 ;
        RECT -18.300 10.020 -17.840 10.200 ;
        RECT -17.510 10.020 -17.050 10.200 ;
        RECT -16.720 10.020 -16.260 10.200 ;
        RECT -15.930 10.020 -15.470 10.200 ;
        RECT -15.140 10.020 -14.680 10.200 ;
        RECT -14.350 10.020 -13.890 10.200 ;
        RECT -13.560 10.020 -13.100 10.200 ;
        RECT -12.770 10.020 -12.310 10.200 ;
        RECT -11.980 10.020 -11.520 10.200 ;
        RECT -11.190 10.020 -10.730 10.200 ;
        RECT -10.400 10.020 -9.940 10.200 ;
        RECT -9.610 10.020 -9.150 10.200 ;
        RECT -8.820 10.020 -8.360 10.200 ;
        RECT -8.030 10.020 -7.570 10.200 ;
        RECT -7.240 10.020 -6.780 10.200 ;
        RECT -6.450 10.020 -5.990 10.200 ;
        RECT -5.660 10.020 -5.200 10.200 ;
        RECT -4.870 10.020 -4.410 10.200 ;
        RECT -4.080 10.020 -3.620 10.200 ;
        RECT -3.290 10.020 -2.830 10.200 ;
        RECT -2.500 10.020 -2.040 10.200 ;
        RECT -1.710 10.020 -1.250 10.200 ;
        RECT -0.920 10.020 -0.460 10.200 ;
        RECT -0.130 10.020 0.330 10.200 ;
        RECT 0.660 10.020 1.120 10.200 ;
        RECT 1.450 10.020 1.910 10.200 ;
        RECT 2.240 10.020 2.700 10.200 ;
        RECT 3.030 10.020 3.490 10.200 ;
        RECT 3.820 10.020 4.280 10.200 ;
        RECT 4.610 10.020 5.070 10.200 ;
        RECT 5.400 10.020 5.860 10.200 ;
        RECT 6.190 10.020 6.650 10.200 ;
        RECT 6.980 10.020 7.440 10.200 ;
        RECT 7.770 10.020 8.230 10.200 ;
        RECT 8.560 10.020 9.020 10.200 ;
        RECT 9.350 10.020 9.810 10.200 ;
        RECT 10.140 10.020 10.600 10.200 ;
        RECT 10.930 10.020 11.390 10.200 ;
        RECT -19.880 8.565 -19.420 8.610 ;
        RECT -19.090 8.565 -18.630 8.610 ;
        RECT -18.300 8.565 -17.840 8.610 ;
        RECT -17.510 8.565 -17.050 8.610 ;
        RECT -16.720 8.565 -16.260 8.610 ;
        RECT -15.930 8.565 -15.470 8.610 ;
        RECT -15.140 8.565 -14.680 8.610 ;
        RECT -14.350 8.565 -13.890 8.610 ;
        RECT -13.560 8.565 -13.100 8.610 ;
        RECT -12.770 8.565 -12.310 8.610 ;
        RECT -11.980 8.565 -11.520 8.610 ;
        RECT -11.190 8.565 -10.730 8.610 ;
        RECT -10.400 8.565 -9.940 8.610 ;
        RECT -9.610 8.565 -9.150 8.610 ;
        RECT -8.820 8.565 -8.360 8.610 ;
        RECT -8.030 8.565 -7.570 8.610 ;
        RECT -7.240 8.565 -6.780 8.610 ;
        RECT -6.450 8.565 -5.990 8.610 ;
        RECT -5.660 8.565 -5.200 8.610 ;
        RECT -4.870 8.565 -4.410 8.610 ;
        RECT -4.080 8.565 -3.620 8.610 ;
        RECT -3.290 8.565 -2.830 8.610 ;
        RECT -2.500 8.565 -2.040 8.610 ;
        RECT -1.710 8.565 -1.250 8.610 ;
        RECT -0.920 8.565 -0.460 8.610 ;
        RECT -0.130 8.565 0.330 8.610 ;
        RECT 0.660 8.565 1.120 8.610 ;
        RECT 1.450 8.565 1.910 8.610 ;
        RECT 2.240 8.565 2.700 8.610 ;
        RECT 3.030 8.565 3.490 8.610 ;
        RECT 3.820 8.565 4.280 8.610 ;
        RECT 4.610 8.565 5.070 8.610 ;
        RECT 5.400 8.565 5.860 8.610 ;
        RECT 6.190 8.565 6.650 8.610 ;
        RECT 6.980 8.565 7.440 8.610 ;
        RECT 7.770 8.565 8.230 8.610 ;
        RECT 8.560 8.565 9.020 8.610 ;
        RECT 9.350 8.565 9.810 8.610 ;
        RECT 10.140 8.565 10.600 8.610 ;
        RECT 10.930 8.565 11.390 8.610 ;
        RECT 12.060 8.565 12.380 10.200 ;
        RECT -20.870 8.245 12.380 8.565 ;
        RECT -21.455 7.595 -18.170 7.915 ;
        RECT 12.060 7.845 12.380 8.245 ;
        RECT -18.490 2.455 -18.170 7.595 ;
        RECT 9.555 7.530 12.380 7.845 ;
        RECT 9.555 7.525 12.060 7.530 ;
        RECT -13.730 4.370 -11.930 4.555 ;
        RECT -13.730 4.200 -13.485 4.370 ;
        RECT -15.565 3.200 -15.190 4.200 ;
        RECT -13.840 3.200 -13.485 4.200 ;
        RECT -15.565 2.980 -15.320 3.200 ;
        RECT -15.140 2.980 -14.680 2.995 ;
        RECT -14.350 2.980 -13.890 2.995 ;
        RECT -13.730 2.980 -13.485 3.200 ;
        RECT -15.565 2.800 -13.485 2.980 ;
        RECT -15.565 2.530 -15.320 2.800 ;
        RECT -15.140 2.765 -14.680 2.800 ;
        RECT -14.350 2.765 -13.890 2.800 ;
        RECT -13.730 2.530 -13.485 2.800 ;
        RECT -12.645 3.200 -12.270 4.200 ;
        RECT -12.645 2.535 -12.400 3.200 ;
        RECT -12.115 2.995 -11.930 4.370 ;
        RECT -7.890 4.390 -6.100 4.575 ;
        RECT -7.890 4.200 -7.645 4.390 ;
        RECT -10.920 3.200 -10.550 4.200 ;
        RECT -12.220 2.975 -11.760 2.995 ;
        RECT -11.430 2.975 -10.970 2.995 ;
        RECT -12.220 2.795 -10.970 2.975 ;
        RECT -12.220 2.765 -11.760 2.795 ;
        RECT -11.430 2.765 -10.970 2.795 ;
        RECT -10.795 2.535 -10.550 3.200 ;
        RECT -18.490 2.180 -16.310 2.455 ;
        RECT -15.565 2.120 -13.485 2.530 ;
        RECT -15.565 2.115 -13.505 2.120 ;
        RECT -15.140 -0.285 -14.685 2.115 ;
        RECT -12.975 2.105 -10.550 2.535 ;
        RECT -9.730 3.200 -9.350 4.200 ;
        RECT -8.000 3.200 -7.645 4.200 ;
        RECT -9.730 2.975 -9.485 3.200 ;
        RECT -9.300 2.975 -8.840 2.995 ;
        RECT -8.510 2.975 -8.050 2.995 ;
        RECT -7.890 2.975 -7.645 3.200 ;
        RECT -9.730 2.795 -7.645 2.975 ;
        RECT -9.730 2.520 -9.485 2.795 ;
        RECT -9.300 2.765 -8.840 2.795 ;
        RECT -8.510 2.765 -8.050 2.795 ;
        RECT -7.890 2.520 -7.645 2.795 ;
        RECT -9.730 2.115 -7.645 2.520 ;
        RECT -6.780 3.200 -6.430 4.200 ;
        RECT -6.780 2.520 -6.535 3.200 ;
        RECT -6.285 2.995 -6.100 4.390 ;
        RECT -5.080 3.200 -4.735 4.200 ;
        RECT -6.380 2.975 -5.920 2.995 ;
        RECT -5.590 2.975 -5.130 2.995 ;
        RECT -6.380 2.795 -5.130 2.975 ;
        RECT -6.380 2.765 -5.920 2.795 ;
        RECT -5.590 2.765 -5.130 2.795 ;
        RECT -4.980 2.520 -4.735 3.200 ;
        RECT -12.975 -0.285 -12.525 2.105 ;
        RECT -11.420 0.105 -10.960 0.430 ;
        RECT -11.420 0.100 -10.955 0.105 ;
        RECT -11.415 -0.125 -10.955 0.100 ;
        RECT -16.035 -0.300 -15.805 -0.285 ;
        RECT -16.105 -1.280 -15.780 -0.300 ;
        RECT -15.245 -1.265 -14.685 -0.285 ;
        RECT -13.865 -0.300 -13.635 -0.285 ;
        RECT -16.035 -1.285 -15.805 -1.280 ;
        RECT -15.245 -1.285 -15.015 -1.265 ;
        RECT -13.940 -1.280 -13.615 -0.300 ;
        RECT -13.075 -1.280 -12.525 -0.285 ;
        RECT -13.865 -1.285 -13.635 -1.280 ;
        RECT -13.075 -1.285 -12.845 -1.280 ;
        RECT -11.280 -1.445 -11.070 -0.125 ;
        RECT -8.620 -0.285 -8.195 2.115 ;
        RECT -6.780 2.110 -4.735 2.520 ;
        RECT -3.895 3.200 -3.510 4.200 ;
        RECT -6.450 -0.285 -5.995 2.110 ;
        RECT -3.895 0.765 -3.665 3.200 ;
        RECT -3.110 3.190 -2.550 4.240 ;
        RECT -2.160 3.200 -1.820 4.200 ;
        RECT -2.050 0.765 -1.820 3.200 ;
        RECT -4.905 -0.125 -4.445 0.430 ;
        RECT -3.895 0.270 -1.820 0.765 ;
        RECT -0.955 3.200 -0.590 4.200 ;
        RECT -0.955 0.760 -0.725 3.200 ;
        RECT -0.180 3.185 0.380 4.235 ;
        RECT 0.760 3.200 1.155 4.200 ;
        RECT 0.925 0.760 1.155 3.200 ;
        RECT 1.940 3.180 2.500 4.230 ;
        RECT 3.535 3.195 4.095 4.245 ;
        RECT 5.840 4.200 6.010 4.220 ;
        RECT 5.810 3.200 6.040 4.200 ;
        RECT 5.840 2.995 6.010 3.200 ;
        RECT 2.380 2.990 2.840 2.995 ;
        RECT 3.170 2.990 3.630 2.995 ;
        RECT 5.295 2.990 6.010 2.995 ;
        RECT 2.380 2.775 6.010 2.990 ;
        RECT 2.380 2.765 2.840 2.775 ;
        RECT 3.170 2.765 3.630 2.775 ;
        RECT 5.295 2.755 6.010 2.775 ;
        RECT -10.905 -0.300 -10.675 -0.285 ;
        RECT -9.525 -0.300 -9.295 -0.285 ;
        RECT -10.915 -1.280 -10.590 -0.300 ;
        RECT -9.580 -1.280 -9.255 -0.300 ;
        RECT -8.735 -1.265 -8.195 -0.285 ;
        RECT -7.355 -0.300 -7.125 -0.285 ;
        RECT -10.905 -1.285 -10.675 -1.280 ;
        RECT -9.525 -1.285 -9.295 -1.280 ;
        RECT -8.735 -1.285 -8.505 -1.265 ;
        RECT -7.425 -1.280 -7.100 -0.300 ;
        RECT -6.565 -1.280 -5.995 -0.285 ;
        RECT -7.355 -1.285 -7.125 -1.280 ;
        RECT -6.565 -1.285 -6.335 -1.280 ;
        RECT -4.775 -1.445 -4.565 -0.125 ;
        RECT -3.425 -0.285 -2.900 0.270 ;
        RECT -0.955 0.255 1.155 0.760 ;
        RECT -2.735 0.065 -2.275 0.105 ;
        RECT -0.565 0.065 -0.105 0.105 ;
        RECT 0.050 0.065 0.610 0.255 ;
        RECT -2.735 -0.105 0.610 0.065 ;
        RECT -2.735 -0.125 -2.275 -0.105 ;
        RECT -0.565 -0.125 -0.105 -0.105 ;
        RECT -4.395 -0.300 -4.165 -0.285 ;
        RECT -4.405 -1.280 -4.080 -0.300 ;
        RECT -4.395 -1.285 -4.165 -1.280 ;
        RECT -3.425 -1.285 -2.785 -0.285 ;
        RECT -11.415 -1.675 -10.955 -1.445 ;
        RECT -4.905 -1.675 -4.445 -1.445 ;
        RECT -3.425 -2.040 -2.900 -1.285 ;
        RECT -2.615 -1.445 -2.420 -0.125 ;
        RECT -0.435 -1.445 -0.240 -0.125 ;
        RECT 0.050 -0.285 0.610 -0.105 ;
        RECT 1.600 0.080 2.060 0.100 ;
        RECT 2.390 0.080 2.850 0.100 ;
        RECT 3.180 0.080 3.640 0.100 ;
        RECT 3.970 0.080 4.430 0.100 ;
        RECT 1.600 -0.095 5.570 0.080 ;
        RECT 1.600 -0.130 2.060 -0.095 ;
        RECT 2.390 -0.130 2.850 -0.095 ;
        RECT 3.180 -0.130 3.640 -0.095 ;
        RECT 3.970 -0.130 4.430 -0.095 ;
        RECT -0.055 -1.285 0.610 -0.285 ;
        RECT 2.010 -1.205 2.420 -0.285 ;
        RECT 3.595 -1.200 4.005 -0.280 ;
        RECT 2.110 -1.290 2.340 -1.205 ;
        RECT 3.690 -1.290 3.920 -1.200 ;
        RECT -2.735 -1.675 -2.275 -1.445 ;
        RECT -0.565 -1.675 -0.105 -1.445 ;
        RECT 1.600 -1.510 2.060 -1.450 ;
        RECT 2.390 -1.510 2.850 -1.450 ;
        RECT 3.180 -1.510 3.640 -1.450 ;
        RECT 3.970 -1.510 4.430 -1.450 ;
        RECT 5.140 -1.510 5.570 -0.095 ;
        RECT 5.795 -0.285 5.985 2.755 ;
        RECT 9.555 2.445 9.875 7.525 ;
        RECT 8.580 2.170 9.875 2.445 ;
        RECT 6.145 0.075 6.605 0.105 ;
        RECT 7.290 0.075 7.645 0.390 ;
        RECT 6.145 -0.075 7.645 0.075 ;
        RECT 6.145 -0.125 6.605 -0.075 ;
        RECT 5.795 -1.285 6.095 -0.285 ;
        RECT 7.290 -0.615 7.645 -0.075 ;
        RECT 8.950 -0.285 9.205 -0.270 ;
        RECT 8.040 -0.615 8.270 -0.285 ;
        RECT 7.290 -0.930 8.270 -0.615 ;
        RECT 6.145 -1.510 6.605 -1.445 ;
        RECT 7.290 -1.510 7.645 -0.930 ;
        RECT 8.040 -1.285 8.270 -0.930 ;
        RECT 8.830 -1.285 9.205 -0.285 ;
        RECT 1.600 -1.660 7.645 -1.510 ;
        RECT 1.600 -1.680 2.060 -1.660 ;
        RECT 2.390 -1.680 2.850 -1.660 ;
        RECT 3.180 -1.680 3.640 -1.660 ;
        RECT 3.970 -1.680 4.430 -1.660 ;
        RECT 6.145 -1.675 6.605 -1.660 ;
        RECT 8.950 -1.835 9.205 -1.285 ;
        RECT -19.545 -2.345 -18.510 -2.040 ;
        RECT -3.600 -2.345 -2.755 -2.040 ;
        RECT 8.950 -2.185 12.945 -1.835 ;
        RECT -19.460 -3.105 -19.125 -2.345 ;
        RECT -20.980 -3.440 -19.125 -3.105 ;
        RECT -20.980 -3.780 -20.645 -3.440 ;
        RECT -20.980 -4.115 12.375 -3.780 ;
        RECT -20.980 -5.625 -20.645 -4.115 ;
        RECT -19.960 -4.210 -19.500 -4.115 ;
        RECT -19.170 -4.210 -18.710 -4.115 ;
        RECT -18.380 -4.210 -17.920 -4.115 ;
        RECT -17.590 -4.210 -17.130 -4.115 ;
        RECT -16.800 -4.210 -16.340 -4.115 ;
        RECT -16.010 -4.210 -15.550 -4.115 ;
        RECT -15.220 -4.210 -14.760 -4.115 ;
        RECT -14.430 -4.210 -13.970 -4.115 ;
        RECT -13.640 -4.210 -13.180 -4.115 ;
        RECT -12.850 -4.210 -12.390 -4.115 ;
        RECT -12.060 -4.210 -11.600 -4.115 ;
        RECT -11.270 -4.210 -10.810 -4.115 ;
        RECT -10.480 -4.210 -10.020 -4.115 ;
        RECT -9.690 -4.210 -9.230 -4.115 ;
        RECT -8.900 -4.210 -8.440 -4.115 ;
        RECT -8.110 -4.210 -7.650 -4.115 ;
        RECT -7.320 -4.210 -6.860 -4.115 ;
        RECT -6.530 -4.210 -6.070 -4.115 ;
        RECT -5.740 -4.210 -5.280 -4.115 ;
        RECT -4.950 -4.210 -4.490 -4.115 ;
        RECT -4.160 -4.210 -3.700 -4.115 ;
        RECT -3.370 -4.210 -2.910 -4.115 ;
        RECT -2.580 -4.210 -2.120 -4.115 ;
        RECT -1.790 -4.210 -1.330 -4.115 ;
        RECT -1.000 -4.210 -0.540 -4.115 ;
        RECT -0.210 -4.210 0.250 -4.115 ;
        RECT 0.580 -4.210 1.040 -4.115 ;
        RECT 1.370 -4.210 1.830 -4.115 ;
        RECT 2.160 -4.210 2.620 -4.115 ;
        RECT 2.950 -4.210 3.410 -4.115 ;
        RECT 3.740 -4.210 4.200 -4.115 ;
        RECT 4.530 -4.210 4.990 -4.115 ;
        RECT 5.320 -4.210 5.780 -4.115 ;
        RECT 6.110 -4.210 6.570 -4.115 ;
        RECT 6.900 -4.210 7.360 -4.115 ;
        RECT 7.690 -4.210 8.150 -4.115 ;
        RECT 8.480 -4.210 8.940 -4.115 ;
        RECT 9.270 -4.210 9.730 -4.115 ;
        RECT 10.060 -4.210 10.520 -4.115 ;
        RECT 10.850 -4.210 11.310 -4.115 ;
        RECT -19.960 -5.625 -19.500 -5.530 ;
        RECT -19.170 -5.625 -18.710 -5.530 ;
        RECT -18.380 -5.625 -17.920 -5.530 ;
        RECT -17.590 -5.625 -17.130 -5.530 ;
        RECT -16.800 -5.625 -16.340 -5.530 ;
        RECT -16.010 -5.625 -15.550 -5.530 ;
        RECT -15.220 -5.625 -14.760 -5.530 ;
        RECT -14.430 -5.625 -13.970 -5.530 ;
        RECT -13.640 -5.625 -13.180 -5.530 ;
        RECT -12.850 -5.625 -12.390 -5.530 ;
        RECT -12.060 -5.625 -11.600 -5.530 ;
        RECT -11.270 -5.625 -10.810 -5.530 ;
        RECT -10.480 -5.625 -10.020 -5.530 ;
        RECT -9.690 -5.625 -9.230 -5.530 ;
        RECT -8.900 -5.625 -8.440 -5.530 ;
        RECT -8.110 -5.625 -7.650 -5.530 ;
        RECT -7.320 -5.625 -6.860 -5.530 ;
        RECT -6.530 -5.625 -6.070 -5.530 ;
        RECT -5.740 -5.625 -5.280 -5.530 ;
        RECT -4.950 -5.625 -4.490 -5.530 ;
        RECT -4.160 -5.625 -3.700 -5.530 ;
        RECT -3.370 -5.625 -2.910 -5.530 ;
        RECT -2.580 -5.625 -2.120 -5.530 ;
        RECT -1.790 -5.625 -1.330 -5.530 ;
        RECT -1.000 -5.625 -0.540 -5.530 ;
        RECT -0.210 -5.625 0.250 -5.530 ;
        RECT 0.580 -5.625 1.040 -5.530 ;
        RECT 1.370 -5.625 1.830 -5.530 ;
        RECT 2.160 -5.625 2.620 -5.530 ;
        RECT 2.950 -5.625 3.410 -5.530 ;
        RECT 3.740 -5.625 4.200 -5.530 ;
        RECT 4.530 -5.625 4.990 -5.530 ;
        RECT 5.320 -5.625 5.780 -5.530 ;
        RECT 6.110 -5.625 6.570 -5.530 ;
        RECT 6.900 -5.625 7.360 -5.530 ;
        RECT 7.690 -5.625 8.150 -5.530 ;
        RECT 8.480 -5.625 8.940 -5.530 ;
        RECT 9.270 -5.625 9.730 -5.530 ;
        RECT 10.060 -5.625 10.520 -5.530 ;
        RECT 10.850 -5.625 11.310 -5.530 ;
        RECT 12.040 -5.625 12.375 -4.115 ;
        RECT -20.980 -6.200 12.375 -5.625 ;
        RECT -20.980 -7.730 -20.645 -6.200 ;
        RECT -19.960 -6.300 -19.500 -6.200 ;
        RECT -19.170 -6.300 -18.710 -6.200 ;
        RECT -18.380 -6.300 -17.920 -6.200 ;
        RECT -17.590 -6.300 -17.130 -6.200 ;
        RECT -16.800 -6.300 -16.340 -6.200 ;
        RECT -16.010 -6.300 -15.550 -6.200 ;
        RECT -15.220 -6.300 -14.760 -6.200 ;
        RECT -14.430 -6.300 -13.970 -6.200 ;
        RECT -13.640 -6.300 -13.180 -6.200 ;
        RECT -12.850 -6.300 -12.390 -6.200 ;
        RECT -12.060 -6.300 -11.600 -6.200 ;
        RECT -11.270 -6.300 -10.810 -6.200 ;
        RECT -10.480 -6.300 -10.020 -6.200 ;
        RECT -9.690 -6.300 -9.230 -6.200 ;
        RECT -8.900 -6.300 -8.440 -6.200 ;
        RECT -8.110 -6.300 -7.650 -6.200 ;
        RECT -7.320 -6.300 -6.860 -6.200 ;
        RECT -6.530 -6.300 -6.070 -6.200 ;
        RECT -5.740 -6.300 -5.280 -6.200 ;
        RECT -4.950 -6.300 -4.490 -6.200 ;
        RECT -4.160 -6.300 -3.700 -6.200 ;
        RECT -3.370 -6.300 -2.910 -6.200 ;
        RECT -2.580 -6.300 -2.120 -6.200 ;
        RECT -1.790 -6.300 -1.330 -6.200 ;
        RECT -1.000 -6.300 -0.540 -6.200 ;
        RECT -0.210 -6.300 0.250 -6.200 ;
        RECT 0.580 -6.300 1.040 -6.200 ;
        RECT 1.370 -6.300 1.830 -6.200 ;
        RECT 2.160 -6.300 2.620 -6.200 ;
        RECT 2.950 -6.300 3.410 -6.200 ;
        RECT 3.740 -6.300 4.200 -6.200 ;
        RECT 4.530 -6.300 4.990 -6.200 ;
        RECT 5.320 -6.300 5.780 -6.200 ;
        RECT 6.110 -6.300 6.570 -6.200 ;
        RECT 6.900 -6.300 7.360 -6.200 ;
        RECT 7.690 -6.300 8.150 -6.200 ;
        RECT 8.480 -6.300 8.940 -6.200 ;
        RECT 9.270 -6.300 9.730 -6.200 ;
        RECT 10.060 -6.300 10.520 -6.200 ;
        RECT 10.850 -6.300 11.310 -6.200 ;
        RECT -19.960 -7.730 -19.500 -7.620 ;
        RECT -19.170 -7.730 -18.710 -7.620 ;
        RECT -18.380 -7.730 -17.920 -7.620 ;
        RECT -17.590 -7.730 -17.130 -7.620 ;
        RECT -16.800 -7.730 -16.340 -7.620 ;
        RECT -16.010 -7.730 -15.550 -7.620 ;
        RECT -15.220 -7.730 -14.760 -7.620 ;
        RECT -14.430 -7.730 -13.970 -7.620 ;
        RECT -13.640 -7.730 -13.180 -7.620 ;
        RECT -12.850 -7.730 -12.390 -7.620 ;
        RECT -12.060 -7.730 -11.600 -7.620 ;
        RECT -11.270 -7.730 -10.810 -7.620 ;
        RECT -10.480 -7.730 -10.020 -7.620 ;
        RECT -9.690 -7.730 -9.230 -7.620 ;
        RECT -8.900 -7.730 -8.440 -7.620 ;
        RECT -8.110 -7.730 -7.650 -7.620 ;
        RECT -7.320 -7.730 -6.860 -7.620 ;
        RECT -6.530 -7.730 -6.070 -7.620 ;
        RECT -5.740 -7.730 -5.280 -7.620 ;
        RECT -4.950 -7.730 -4.490 -7.620 ;
        RECT -4.160 -7.730 -3.700 -7.620 ;
        RECT -3.370 -7.730 -2.910 -7.620 ;
        RECT -2.580 -7.730 -2.120 -7.620 ;
        RECT -1.790 -7.730 -1.330 -7.620 ;
        RECT -1.000 -7.730 -0.540 -7.620 ;
        RECT -0.210 -7.730 0.250 -7.620 ;
        RECT 0.580 -7.730 1.040 -7.620 ;
        RECT 1.370 -7.730 1.830 -7.620 ;
        RECT 2.160 -7.730 2.620 -7.620 ;
        RECT 2.950 -7.730 3.410 -7.620 ;
        RECT 3.740 -7.730 4.200 -7.620 ;
        RECT 4.530 -7.730 4.990 -7.620 ;
        RECT 5.320 -7.730 5.780 -7.620 ;
        RECT 6.110 -7.730 6.570 -7.620 ;
        RECT 6.900 -7.730 7.360 -7.620 ;
        RECT 7.690 -7.730 8.150 -7.620 ;
        RECT 8.480 -7.730 8.940 -7.620 ;
        RECT 9.270 -7.730 9.730 -7.620 ;
        RECT 10.060 -7.730 10.520 -7.620 ;
        RECT 10.850 -7.730 11.310 -7.620 ;
        RECT 12.040 -7.730 12.375 -6.200 ;
        RECT -20.980 -8.305 12.375 -7.730 ;
        RECT -20.980 -9.780 -20.645 -8.305 ;
        RECT -19.960 -8.390 -19.500 -8.305 ;
        RECT -19.170 -8.390 -18.710 -8.305 ;
        RECT -18.380 -8.390 -17.920 -8.305 ;
        RECT -17.590 -8.390 -17.130 -8.305 ;
        RECT -16.800 -8.390 -16.340 -8.305 ;
        RECT -16.010 -8.390 -15.550 -8.305 ;
        RECT -15.220 -8.390 -14.760 -8.305 ;
        RECT -14.430 -8.390 -13.970 -8.305 ;
        RECT -13.640 -8.390 -13.180 -8.305 ;
        RECT -12.850 -8.390 -12.390 -8.305 ;
        RECT -12.060 -8.390 -11.600 -8.305 ;
        RECT -11.270 -8.390 -10.810 -8.305 ;
        RECT -10.480 -8.390 -10.020 -8.305 ;
        RECT -9.690 -8.390 -9.230 -8.305 ;
        RECT -8.900 -8.390 -8.440 -8.305 ;
        RECT -8.110 -8.390 -7.650 -8.305 ;
        RECT -7.320 -8.390 -6.860 -8.305 ;
        RECT -6.530 -8.390 -6.070 -8.305 ;
        RECT -5.740 -8.390 -5.280 -8.305 ;
        RECT -4.950 -8.390 -4.490 -8.305 ;
        RECT -4.160 -8.390 -3.700 -8.305 ;
        RECT -3.370 -8.390 -2.910 -8.305 ;
        RECT -2.580 -8.390 -2.120 -8.305 ;
        RECT -1.790 -8.390 -1.330 -8.305 ;
        RECT -1.000 -8.390 -0.540 -8.305 ;
        RECT -0.210 -8.390 0.250 -8.305 ;
        RECT 0.580 -8.390 1.040 -8.305 ;
        RECT 1.370 -8.390 1.830 -8.305 ;
        RECT 2.160 -8.390 2.620 -8.305 ;
        RECT 2.950 -8.390 3.410 -8.305 ;
        RECT 3.740 -8.390 4.200 -8.305 ;
        RECT 4.530 -8.390 4.990 -8.305 ;
        RECT 5.320 -8.390 5.780 -8.305 ;
        RECT 6.110 -8.390 6.570 -8.305 ;
        RECT 6.900 -8.390 7.360 -8.305 ;
        RECT 7.690 -8.390 8.150 -8.305 ;
        RECT 8.480 -8.390 8.940 -8.305 ;
        RECT 9.270 -8.390 9.730 -8.305 ;
        RECT 10.060 -8.390 10.520 -8.305 ;
        RECT 10.850 -8.390 11.310 -8.305 ;
        RECT -19.960 -9.780 -19.500 -9.710 ;
        RECT -19.170 -9.780 -18.710 -9.710 ;
        RECT -18.380 -9.780 -17.920 -9.710 ;
        RECT -17.590 -9.780 -17.130 -9.710 ;
        RECT -16.800 -9.780 -16.340 -9.710 ;
        RECT -16.010 -9.780 -15.550 -9.710 ;
        RECT -15.220 -9.780 -14.760 -9.710 ;
        RECT -14.430 -9.780 -13.970 -9.710 ;
        RECT -13.640 -9.780 -13.180 -9.710 ;
        RECT -12.850 -9.780 -12.390 -9.710 ;
        RECT -12.060 -9.780 -11.600 -9.710 ;
        RECT -11.270 -9.780 -10.810 -9.710 ;
        RECT -10.480 -9.780 -10.020 -9.710 ;
        RECT -9.690 -9.780 -9.230 -9.710 ;
        RECT -8.900 -9.780 -8.440 -9.710 ;
        RECT -8.110 -9.780 -7.650 -9.710 ;
        RECT -7.320 -9.780 -6.860 -9.710 ;
        RECT -6.530 -9.780 -6.070 -9.710 ;
        RECT -5.740 -9.780 -5.280 -9.710 ;
        RECT -4.950 -9.780 -4.490 -9.710 ;
        RECT -4.160 -9.780 -3.700 -9.710 ;
        RECT -3.370 -9.780 -2.910 -9.710 ;
        RECT -2.580 -9.780 -2.120 -9.710 ;
        RECT -1.790 -9.780 -1.330 -9.710 ;
        RECT -1.000 -9.780 -0.540 -9.710 ;
        RECT -0.210 -9.780 0.250 -9.710 ;
        RECT 0.580 -9.780 1.040 -9.710 ;
        RECT 1.370 -9.780 1.830 -9.710 ;
        RECT 2.160 -9.780 2.620 -9.710 ;
        RECT 2.950 -9.780 3.410 -9.710 ;
        RECT 3.740 -9.780 4.200 -9.710 ;
        RECT 4.530 -9.780 4.990 -9.710 ;
        RECT 5.320 -9.780 5.780 -9.710 ;
        RECT 6.110 -9.780 6.570 -9.710 ;
        RECT 6.900 -9.780 7.360 -9.710 ;
        RECT 7.690 -9.780 8.150 -9.710 ;
        RECT 8.480 -9.780 8.940 -9.710 ;
        RECT 9.270 -9.780 9.730 -9.710 ;
        RECT 10.060 -9.780 10.520 -9.710 ;
        RECT 10.850 -9.780 11.310 -9.710 ;
        RECT 12.040 -9.780 12.375 -8.305 ;
        RECT -20.980 -10.115 12.375 -9.780 ;
        RECT 12.595 -11.820 12.945 -2.185 ;
        RECT -19.080 -12.130 -16.975 -11.880 ;
        RECT -18.960 -13.470 -17.170 -12.130 ;
        RECT 8.020 -12.170 12.945 -11.820 ;
        RECT -19.080 -13.720 -16.975 -13.470 ;
        RECT 8.075 -13.720 10.180 -13.470 ;
        RECT 8.105 -15.060 9.895 -13.720 ;
        RECT -19.080 -15.310 -16.975 -15.060 ;
        RECT 8.075 -15.310 10.180 -15.060 ;
        RECT -18.960 -16.650 -17.170 -15.310 ;
        RECT -19.080 -16.900 -16.975 -16.650 ;
      LAYER met2 ;
        RECT -3.915 3.185 4.105 4.235 ;
        RECT -17.225 2.180 -10.485 2.455 ;
        RECT -6.885 2.170 9.875 2.445 ;
        RECT -11.465 0.350 -10.930 0.400 ;
        RECT -4.935 0.350 -4.415 0.400 ;
        RECT 7.290 0.350 7.645 0.390 ;
        RECT -11.465 0.140 7.645 0.350 ;
        RECT -16.105 -1.280 -10.590 -0.300 ;
        RECT -9.580 -1.280 -4.080 -0.300 ;
        RECT 1.985 -1.215 2.425 0.140 ;
        RECT 3.585 -1.215 4.025 0.140 ;
        RECT 5.140 -1.650 5.575 0.140 ;
        RECT 7.290 -1.685 7.645 0.140 ;
        RECT -19.545 -2.345 -2.755 -2.040 ;
  END
END sky130_ef_ip__opamp
END LIBRARY

