magic
tech sky130A
magscale 1 2
timestamp 1723064828
<< error_s >>
rect 111 -1798 157 -1772
rect 83 -1826 185 -1800
rect 596 -2029 613 -1413
rect 650 -2078 667 -1462
rect 1177 -1474 1292 -1462
rect 1184 -1508 1292 -1474
rect 1177 -1520 1292 -1508
rect 1234 -1575 1292 -1520
rect 1275 -2124 1292 -1575
rect 1293 -1575 1358 -1539
rect 1293 -1633 1444 -1575
rect 1293 -2124 1387 -1633
rect 1293 -2190 1358 -2124
rect 1766 -2219 1813 -1586
rect 1820 -2273 1867 -1640
rect 2763 -2272 2766 -1652
rect 2797 -2284 2831 -1586
rect 3093 -1674 3127 -1588
rect 3068 -1740 3163 -1674
rect 3068 -1798 3279 -1740
rect 34945 -1752 35060 -1740
rect 34952 -1786 35060 -1752
rect 34945 -1798 35060 -1786
rect 2797 -2303 2800 -2284
rect 3068 -2337 3192 -1798
rect 35002 -1853 35060 -1798
rect 3268 -2171 3279 -1971
rect 3068 -2373 3163 -2337
rect 35043 -2402 35060 -1853
rect 35061 -1853 35126 -1817
rect 35061 -1911 35212 -1853
rect 35061 -2402 35155 -1911
rect 35061 -2468 35126 -2402
rect 54336 -2497 54383 -1864
rect 54815 -1918 54910 -1899
rect 54390 -2551 54437 -1918
rect 54729 -1965 54910 -1918
rect 54815 -2023 55026 -1965
rect 54815 -2562 54939 -2023
rect 55015 -2396 55026 -2196
rect 54815 -2598 54928 -2562
rect 54881 -2616 54928 -2598
rect 55348 -2627 55365 -2011
rect 55402 -2676 55419 -2060
rect 56027 -2722 56044 -2106
rect 56081 -2771 56098 -2155
rect 56706 -2817 56723 -2201
rect 56760 -2866 56777 -2250
rect 57287 -2262 57402 -2250
rect 57294 -2296 57402 -2262
rect 57287 -2308 57402 -2296
rect 57344 -2363 57402 -2308
rect 57385 -2912 57402 -2363
rect 57403 -2363 57468 -2327
rect 57403 -2421 57554 -2363
rect 57403 -2912 57497 -2421
rect 57403 -2978 57468 -2912
rect 57876 -3007 57923 -2374
rect 57930 -3061 57977 -2428
rect 58367 -3072 58414 -2439
rect 58421 -3126 58468 -2493
rect 58858 -3137 58905 -2504
rect 59337 -2558 59432 -2539
rect 58912 -3191 58959 -2558
rect 59251 -2605 59432 -2558
rect 59337 -2663 59548 -2605
rect 59337 -3202 59461 -2663
rect 59537 -3036 59548 -2836
rect 59337 -3238 59450 -3202
rect 59403 -3256 59450 -3238
rect 60028 -3267 60045 -2651
rect 60082 -3316 60099 -2700
rect 60609 -2712 60724 -2700
rect 60616 -2746 60724 -2712
rect 60609 -2758 60724 -2746
rect 60666 -2813 60724 -2758
rect 60707 -3362 60724 -2813
rect 60725 -2813 60790 -2777
rect 60725 -2871 60876 -2813
rect 60725 -3362 60819 -2871
rect 60725 -3428 60790 -3362
rect 61198 -3457 61245 -2824
rect 61252 -3511 61299 -2878
rect 61689 -3522 61736 -2889
rect 62168 -2943 62263 -2924
rect 61743 -3576 61790 -2943
rect 62082 -2990 62263 -2943
rect 62168 -3048 62379 -2990
rect 62168 -3587 62292 -3048
rect 62368 -3421 62379 -3221
rect 94102 -3441 94160 -3289
rect 94173 -3441 94226 -3405
rect 94173 -3475 94312 -3441
rect 62168 -3623 62281 -3587
rect 62234 -3641 62281 -3623
rect 94173 -3652 94243 -3475
rect 94173 -3718 94226 -3652
rect 94488 -3735 94503 -3441
rect 94510 -3735 94557 -3387
rect 94959 -3559 94994 -3505
rect 94522 -3769 94537 -3735
rect 94979 -3788 94982 -3559
rect 95013 -3593 95048 -3559
rect 95272 -3593 95307 -3559
rect 95013 -3800 95047 -3593
rect 95273 -3612 95307 -3593
rect 95013 -3819 95016 -3800
rect 95292 -3853 95307 -3612
rect 95326 -3646 95361 -3612
rect 95326 -3853 95360 -3646
rect 95326 -3887 95341 -3853
rect 95690 -3885 95714 -3517
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__res_generic_l1_M53S24  R3
timestamp 1723064828
transform 1 0 95673 0 1 -3701
box -17 -241 41 241
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XDD1 ~/Tesis/magic
timestamp 1723064828
transform 1 0 94356 0 1 -3588
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XDD2
timestamp 1723064828
transform 1 0 95160 0 1 -3706
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XDD3
timestamp 1723064828
transform 1 0 95473 0 1 -3759
box -183 -183 183 183
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM1 ~/Tesis/magic
timestamp 1723064828
transform 1 0 58663 0 1 -2815
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM2
timestamp 1723064828
transform 1 0 59154 0 1 -2880
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM3 ~/Tesis/magic
timestamp 1723064828
transform 1 0 59724 0 1 -2936
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM4
timestamp 1723064828
transform 1 0 292 0 1 -1698
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM5
timestamp 1723064828
transform 1 0 971 0 1 -1793
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM6
timestamp 1723064828
transform 1 0 60403 0 1 -3031
box -387 -397 387 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM7
timestamp 1723064828
transform 1 0 61003 0 1 -3135
box -278 -358 278 358
use sky130_fd_pr__nfet_03v3_nvt_UNEQ2N  XM8 ~/Tesis/magic
timestamp 1723064828
transform 1 0 61494 0 1 -3200
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM9
timestamp 1723064828
transform 1 0 1571 0 1 -1897
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_H7BQ24  XM10 ~/Tesis/magic
timestamp 1723064828
transform 1 0 2299 0 1 -1962
box -515 -358 515 358
use sky130_fd_pr__nfet_03v3_nvt_UNEQ2N  XM11
timestamp 1723064828
transform 1 0 61985 0 1 -3265
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_54RBUL  XM12 ~/Tesis/magic
timestamp 1723064828
transform 1 0 78197 0 1 -3321
box -16029 -397 16029 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM13
timestamp 1723064828
transform 1 0 94752 0 1 -3478
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_54RBUL  XM20
timestamp 1723064828
transform 1 0 19097 0 1 -2071
box -16029 -397 16029 397
use sky130_fd_pr__nfet_g5v0d10v5_A3MY9Q  XM22 ~/Tesis/magic
timestamp 1723064828
transform 1 0 44740 0 1 -2175
box -9679 -358 9679 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM24
timestamp 1723064828
transform 1 0 54632 0 1 -2240
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM25 ~/Tesis/magic
timestamp 1723064828
transform 1 0 55123 0 1 -2296
box -308 -397 308 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM26
timestamp 1723064828
transform 1 0 55723 0 1 -2391
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM27
timestamp 1723064828
transform 1 0 56402 0 1 -2486
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM28
timestamp 1723064828
transform 1 0 57081 0 1 -2581
box -387 -397 387 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM29
timestamp 1723064828
transform 1 0 57681 0 1 -2685
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM30
timestamp 1723064828
transform 1 0 58172 0 1 -2750
box -278 -358 278 358
use sky130_fd_pr__res_xhigh_po_0p35_E5287M  XR1 ~/Tesis/magic
timestamp 1723064828
transform 1 0 2962 0 1 8209
box -201 -10582 201 10582
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 128 0 0 0 vss
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 128 0 0 0 out
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 128 0 0 0 inm
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 128 0 0 0 inp
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 128 0 0 0 ena
port 5 nsew
<< end >>
